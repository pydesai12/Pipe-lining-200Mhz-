
module calc_DW01_add_6 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n29, n30, n31,
         n32, n35, n37, n38, n39, n40, n41, n43, n45, n46, n47, n48, n49, n51,
         n53, n54, n55, n56, n57, n59, n61, n62, n63, n64, n65, n67, n69, n70,
         n71, n72, n74, n76, n77, n79, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n167, n174, n180, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n312, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311;

  CFA1X1 U3 ( .A(A[30]), .B(n30), .CI(B[30]), .CO(n29), .S(SUM[30]) );
  CFA1X1 U4 ( .A(A[29]), .B(n31), .CI(B[29]), .CO(n30), .S(SUM[29]) );
  CFA1X1 U5 ( .A(A[28]), .B(n32), .CI(B[28]), .CO(n31), .S(SUM[28]) );
  CFA1X1 U6 ( .A(A[27]), .B(n305), .CI(B[27]), .CO(n32), .S(SUM[27]) );
  COND1X1 U227 ( .A(n39), .B(n41), .C(n40), .Z(n38) );
  CNR2XL U228 ( .A(n160), .B(n157), .Z(n155) );
  CNR2X1 U229 ( .A(B[2]), .B(A[2]), .Z(n160) );
  COND1X1 U230 ( .A(n164), .B(n167), .C(n165), .Z(n163) );
  CNR2X1 U231 ( .A(B[1]), .B(A[1]), .Z(n164) );
  CNR2XL U232 ( .A(B[4]), .B(A[4]), .Z(n151) );
  CND2X1 U233 ( .A(B[4]), .B(A[4]), .Z(n152) );
  CANR1XL U234 ( .A(n79), .B(n304), .C(n74), .Z(n72) );
  COND1XL U235 ( .A(n134), .B(n154), .C(n135), .Z(n133) );
  CANR1X1 U236 ( .A(n307), .B(n70), .C(n67), .Z(n65) );
  CANR1XL U237 ( .A(n311), .B(n46), .C(n43), .Z(n41) );
  CAN2X2 U238 ( .A(n303), .B(n167), .Z(SUM[0]) );
  CND2XL U239 ( .A(n193), .B(n161), .Z(n26) );
  CND2XL U240 ( .A(n190), .B(n147), .Z(n23) );
  CNIVX1 U241 ( .A(n312), .Z(SUM[1]) );
  CND2XL U242 ( .A(B[0]), .B(A[0]), .Z(n167) );
  COND1X1 U243 ( .A(n47), .B(n49), .C(n48), .Z(n46) );
  CND2XL U244 ( .A(B[10]), .B(A[10]), .Z(n121) );
  CNR2XL U245 ( .A(B[10]), .B(A[10]), .Z(n120) );
  CANR1X1 U246 ( .A(n155), .B(n163), .C(n156), .Z(n154) );
  CNR2X1 U247 ( .A(n301), .B(n85), .Z(n83) );
  COND1XL U248 ( .A(n86), .B(n112), .C(n87), .Z(n85) );
  COND1X1 U249 ( .A(n71), .B(n83), .C(n72), .Z(n70) );
  CANR1X1 U250 ( .A(n308), .B(n62), .C(n59), .Z(n57) );
  COND1X1 U251 ( .A(n55), .B(n57), .C(n56), .Z(n300) );
  CAN2X1 U252 ( .A(n133), .B(n84), .Z(n301) );
  CIVXL U253 ( .A(n83), .Z(n82) );
  CNR2X1 U254 ( .A(B[14]), .B(A[14]), .Z(n95) );
  CND2X1 U255 ( .A(B[14]), .B(A[14]), .Z(n96) );
  CND2XL U256 ( .A(B[2]), .B(A[2]), .Z(n161) );
  CANR1X1 U257 ( .A(n309), .B(n300), .C(n51), .Z(n49) );
  CANR1XL U258 ( .A(n145), .B(n136), .C(n137), .Z(n135) );
  CND2XL U259 ( .A(n194), .B(n165), .Z(n27) );
  CNR2X1 U260 ( .A(B[12]), .B(A[12]), .Z(n107) );
  COND1X1 U261 ( .A(n63), .B(n65), .C(n64), .Z(n62) );
  CND2XL U262 ( .A(n144), .B(n136), .Z(n134) );
  CNR2XL U263 ( .A(n141), .B(n138), .Z(n136) );
  CNR2XL U264 ( .A(n107), .B(n102), .Z(n100) );
  CNR2XL U265 ( .A(n130), .B(n127), .Z(n125) );
  CND2IX1 U266 ( .B(n47), .A(n48), .Z(n5) );
  CND2IX1 U267 ( .B(n39), .A(n40), .Z(n3) );
  CNR2XL U268 ( .A(n120), .B(n115), .Z(n113) );
  CEOXL U269 ( .A(n7), .B(n57), .Z(SUM[21]) );
  CND2IX1 U270 ( .B(n63), .A(n64), .Z(n9) );
  CND2XL U271 ( .A(n183), .B(n108), .Z(n16) );
  CND2XL U272 ( .A(n180), .B(n91), .Z(n13) );
  CND2XL U273 ( .A(n185), .B(n121), .Z(n18) );
  CEOXL U274 ( .A(n167), .B(n27), .Z(n312) );
  CND2XL U275 ( .A(n187), .B(n131), .Z(n20) );
  CIVXL U276 ( .A(n151), .Z(n191) );
  CENX1 U277 ( .A(n302), .B(n29), .Z(SUM[31]) );
  CENX1 U278 ( .A(A[31]), .B(B[31]), .Z(n302) );
  CNR2XL U279 ( .A(B[8]), .B(A[8]), .Z(n130) );
  CNR2XL U280 ( .A(B[19]), .B(A[19]), .Z(n63) );
  CNR2XL U281 ( .A(B[21]), .B(A[21]), .Z(n55) );
  CNR2XL U282 ( .A(B[23]), .B(A[23]), .Z(n47) );
  CND2XL U283 ( .A(B[16]), .B(A[16]), .Z(n81) );
  CND2XL U284 ( .A(B[17]), .B(A[17]), .Z(n76) );
  CND2XL U285 ( .A(B[18]), .B(A[18]), .Z(n69) );
  CND2XL U286 ( .A(B[20]), .B(A[20]), .Z(n61) );
  CND2XL U287 ( .A(B[22]), .B(A[22]), .Z(n53) );
  CND2XL U288 ( .A(B[6]), .B(A[6]), .Z(n142) );
  CND2XL U289 ( .A(B[1]), .B(A[1]), .Z(n165) );
  CND2XL U290 ( .A(B[3]), .B(A[3]), .Z(n158) );
  CND2XL U291 ( .A(B[9]), .B(A[9]), .Z(n128) );
  CND2XL U292 ( .A(B[5]), .B(A[5]), .Z(n147) );
  CND2XL U293 ( .A(B[7]), .B(A[7]), .Z(n139) );
  CND2XL U294 ( .A(B[13]), .B(A[13]), .Z(n103) );
  CND2XL U295 ( .A(B[11]), .B(A[11]), .Z(n116) );
  CND2XL U296 ( .A(B[19]), .B(A[19]), .Z(n64) );
  CND2XL U297 ( .A(B[21]), .B(A[21]), .Z(n56) );
  CND2XL U298 ( .A(B[23]), .B(A[23]), .Z(n48) );
  COR2XL U299 ( .A(B[17]), .B(A[17]), .Z(n304) );
  COR2XL U300 ( .A(B[16]), .B(A[16]), .Z(n306) );
  COR2XL U301 ( .A(B[22]), .B(A[22]), .Z(n309) );
  COR2XL U302 ( .A(B[18]), .B(A[18]), .Z(n307) );
  COR2XL U303 ( .A(B[20]), .B(A[20]), .Z(n308) );
  CNR2XL U304 ( .A(B[25]), .B(A[25]), .Z(n39) );
  CND2XL U305 ( .A(B[24]), .B(A[24]), .Z(n45) );
  CND2XL U306 ( .A(B[26]), .B(A[26]), .Z(n37) );
  CND2XL U307 ( .A(B[25]), .B(A[25]), .Z(n40) );
  COR2XL U308 ( .A(B[26]), .B(A[26]), .Z(n310) );
  COR2XL U309 ( .A(B[24]), .B(A[24]), .Z(n311) );
  COR2XL U310 ( .A(B[0]), .B(A[0]), .Z(n303) );
  CNR2X1 U311 ( .A(n111), .B(n86), .Z(n84) );
  CND2X1 U312 ( .A(n100), .B(n88), .Z(n86) );
  CND2X1 U313 ( .A(n125), .B(n113), .Z(n111) );
  COND1XL U314 ( .A(n98), .B(n109), .C(n99), .Z(n97) );
  COND1XL U315 ( .A(n111), .B(n132), .C(n112), .Z(n110) );
  CANR1XL U316 ( .A(n144), .B(n153), .C(n145), .Z(n143) );
  COND1XL U317 ( .A(n123), .B(n132), .C(n124), .Z(n122) );
  COND1XL U318 ( .A(n55), .B(n57), .C(n56), .Z(n54) );
  CND2X1 U319 ( .A(n306), .B(n304), .Z(n71) );
  COND1XL U320 ( .A(n161), .B(n157), .C(n158), .Z(n156) );
  COND1XL U321 ( .A(n108), .B(n102), .C(n103), .Z(n101) );
  COND1XL U322 ( .A(n131), .B(n127), .C(n128), .Z(n126) );
  CANR1XL U323 ( .A(n126), .B(n113), .C(n114), .Z(n112) );
  COND1XL U324 ( .A(n121), .B(n115), .C(n116), .Z(n114) );
  COND1XL U325 ( .A(n152), .B(n146), .C(n147), .Z(n145) );
  CANR1XL U326 ( .A(n101), .B(n88), .C(n89), .Z(n87) );
  COND1XL U327 ( .A(n96), .B(n90), .C(n91), .Z(n89) );
  CNR2X1 U328 ( .A(n95), .B(n90), .Z(n88) );
  COND1XL U329 ( .A(n142), .B(n138), .C(n139), .Z(n137) );
  CNR2X1 U330 ( .A(n151), .B(n146), .Z(n144) );
  CENX1 U331 ( .A(n38), .B(n2), .Z(SUM[26]) );
  CND2X1 U332 ( .A(n310), .B(n37), .Z(n2) );
  CENX1 U333 ( .A(n62), .B(n8), .Z(SUM[20]) );
  CND2X1 U334 ( .A(n308), .B(n61), .Z(n8) );
  CENX1 U335 ( .A(n54), .B(n6), .Z(SUM[22]) );
  CND2X1 U336 ( .A(n309), .B(n53), .Z(n6) );
  CENX1 U337 ( .A(n46), .B(n4), .Z(SUM[24]) );
  CND2X1 U338 ( .A(n311), .B(n45), .Z(n4) );
  CEOX1 U339 ( .A(n13), .B(n92), .Z(SUM[15]) );
  CANR1XL U340 ( .A(n93), .B(n97), .C(n94), .Z(n92) );
  CND2X1 U341 ( .A(n174), .B(n56), .Z(n7) );
  CENX1 U342 ( .A(n159), .B(n25), .Z(SUM[3]) );
  CND2X1 U343 ( .A(n192), .B(n158), .Z(n25) );
  COND1XL U344 ( .A(n160), .B(n162), .C(n161), .Z(n159) );
  CENX1 U345 ( .A(n153), .B(n24), .Z(SUM[4]) );
  CND2X1 U346 ( .A(n191), .B(n152), .Z(n24) );
  CENX1 U347 ( .A(n140), .B(n21), .Z(SUM[7]) );
  CND2X1 U348 ( .A(n188), .B(n139), .Z(n21) );
  COND1XL U349 ( .A(n141), .B(n143), .C(n142), .Z(n140) );
  CENX1 U350 ( .A(n129), .B(n19), .Z(SUM[9]) );
  CND2X1 U351 ( .A(n186), .B(n128), .Z(n19) );
  COND1XL U352 ( .A(n130), .B(n132), .C(n131), .Z(n129) );
  CENX1 U353 ( .A(n122), .B(n18), .Z(SUM[10]) );
  CENX1 U354 ( .A(n97), .B(n14), .Z(SUM[14]) );
  CND2X1 U355 ( .A(n93), .B(n96), .Z(n14) );
  CENX1 U356 ( .A(n82), .B(n12), .Z(SUM[16]) );
  CND2X1 U357 ( .A(n306), .B(n81), .Z(n12) );
  CENX1 U358 ( .A(n70), .B(n10), .Z(SUM[18]) );
  CND2X1 U359 ( .A(n307), .B(n69), .Z(n10) );
  CEOX1 U360 ( .A(n26), .B(n162), .Z(SUM[2]) );
  CEOX1 U361 ( .A(n23), .B(n148), .Z(SUM[5]) );
  CANR1XL U362 ( .A(n191), .B(n153), .C(n150), .Z(n148) );
  CEOX1 U363 ( .A(n22), .B(n143), .Z(SUM[6]) );
  CND2X1 U364 ( .A(n189), .B(n142), .Z(n22) );
  CEOX1 U365 ( .A(n20), .B(n132), .Z(SUM[8]) );
  CEOX1 U366 ( .A(n17), .B(n117), .Z(SUM[11]) );
  CND2X1 U367 ( .A(n184), .B(n116), .Z(n17) );
  CANR1XL U368 ( .A(n185), .B(n122), .C(n119), .Z(n117) );
  CEOX1 U369 ( .A(n16), .B(n109), .Z(SUM[12]) );
  CEOX1 U370 ( .A(n15), .B(n104), .Z(SUM[13]) );
  CND2X1 U371 ( .A(n182), .B(n103), .Z(n15) );
  CANR1XL U372 ( .A(n183), .B(n110), .C(n106), .Z(n104) );
  CEOX1 U373 ( .A(n11), .B(n77), .Z(SUM[17]) );
  CND2X1 U374 ( .A(n304), .B(n76), .Z(n11) );
  CANR1XL U375 ( .A(n306), .B(n82), .C(n79), .Z(n77) );
  CNR2X1 U376 ( .A(B[5]), .B(A[5]), .Z(n146) );
  CNR2X1 U377 ( .A(B[13]), .B(A[13]), .Z(n102) );
  CNR2X1 U378 ( .A(B[7]), .B(A[7]), .Z(n138) );
  CNR2X1 U379 ( .A(B[9]), .B(A[9]), .Z(n127) );
  CNR2X1 U380 ( .A(B[11]), .B(A[11]), .Z(n115) );
  CNR2X1 U381 ( .A(B[3]), .B(A[3]), .Z(n157) );
  CNR2X1 U382 ( .A(B[6]), .B(A[6]), .Z(n141) );
  CNR2X1 U383 ( .A(B[15]), .B(A[15]), .Z(n90) );
  CAOR1X1 U384 ( .A(n310), .B(n38), .C(n35), .Z(n305) );
  CND2X1 U385 ( .A(B[12]), .B(A[12]), .Z(n108) );
  CND2X1 U386 ( .A(B[8]), .B(A[8]), .Z(n131) );
  CEOXL U387 ( .A(n5), .B(n49), .Z(SUM[23]) );
  CEOXL U388 ( .A(n9), .B(n65), .Z(SUM[19]) );
  CEOXL U389 ( .A(n3), .B(n41), .Z(SUM[25]) );
  CND2X1 U390 ( .A(B[15]), .B(A[15]), .Z(n91) );
  CIVX2 U391 ( .A(n101), .Z(n99) );
  CIVX2 U392 ( .A(n100), .Z(n98) );
  CIVX2 U393 ( .A(n96), .Z(n94) );
  CIVX2 U394 ( .A(n81), .Z(n79) );
  CIVX2 U395 ( .A(n76), .Z(n74) );
  CIVX2 U396 ( .A(n69), .Z(n67) );
  CIVX2 U397 ( .A(n61), .Z(n59) );
  CIVX2 U398 ( .A(n53), .Z(n51) );
  CIVX2 U399 ( .A(n45), .Z(n43) );
  CIVX2 U400 ( .A(n37), .Z(n35) );
  CIVX2 U401 ( .A(n164), .Z(n194) );
  CIVX2 U402 ( .A(n160), .Z(n193) );
  CIVX2 U403 ( .A(n157), .Z(n192) );
  CIVX2 U404 ( .A(n146), .Z(n190) );
  CIVX2 U405 ( .A(n141), .Z(n189) );
  CIVX2 U406 ( .A(n138), .Z(n188) );
  CIVX2 U407 ( .A(n130), .Z(n187) );
  CIVX2 U408 ( .A(n127), .Z(n186) );
  CIVX2 U409 ( .A(n115), .Z(n184) );
  CIVX2 U410 ( .A(n102), .Z(n182) );
  CIVX2 U411 ( .A(n95), .Z(n93) );
  CIVX2 U412 ( .A(n90), .Z(n180) );
  CIVX2 U413 ( .A(n55), .Z(n174) );
  CIVX2 U414 ( .A(n163), .Z(n162) );
  CIVX2 U415 ( .A(n154), .Z(n153) );
  CIVX2 U416 ( .A(n152), .Z(n150) );
  CIVX2 U417 ( .A(n133), .Z(n132) );
  CIVX2 U418 ( .A(n126), .Z(n124) );
  CIVX2 U419 ( .A(n125), .Z(n123) );
  CIVX2 U420 ( .A(n121), .Z(n119) );
  CIVX2 U421 ( .A(n120), .Z(n185) );
  CIVX2 U422 ( .A(n110), .Z(n109) );
  CIVX2 U423 ( .A(n108), .Z(n106) );
  CIVX2 U424 ( .A(n107), .Z(n183) );
endmodule


module calc_DW01_add_7 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n30, n31,
         n32, n35, n37, n38, n39, n40, n41, n43, n45, n46, n47, n48, n49, n51,
         n53, n54, n55, n56, n57, n59, n61, n62, n63, n64, n65, n67, n69, n70,
         n71, n72, n73, n75, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n165, n176, n178, n179, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n308, n299, n300, n301, n302, n303, n304, n305, n306, n307;

  CFA1X1 U3 ( .A(B[30]), .B(n31), .CI(A[30]), .CO(n30), .S(SUM[30]) );
  CFA1X1 U4 ( .A(B[29]), .B(n32), .CI(A[29]), .CO(n31), .S(SUM[29]) );
  CFA1X1 U5 ( .A(B[28]), .B(n301), .CI(A[28]), .CO(n32), .S(SUM[28]) );
  COND1X1 U58 ( .A(n63), .B(n65), .C(n64), .Z(n62) );
  CENXL U227 ( .A(n78), .B(n12), .Z(SUM[17]) );
  CANR1X1 U228 ( .A(n302), .B(n78), .C(n75), .Z(n73) );
  COND1X1 U229 ( .A(n79), .B(n81), .C(n80), .Z(n78) );
  CENXL U230 ( .A(n70), .B(n10), .Z(SUM[19]) );
  CANR1X1 U231 ( .A(n304), .B(n70), .C(n67), .Z(n65) );
  COND1X1 U232 ( .A(n71), .B(n73), .C(n72), .Z(n70) );
  COND1X2 U233 ( .A(n39), .B(n41), .C(n40), .Z(n38) );
  CANR1X2 U234 ( .A(n307), .B(n46), .C(n43), .Z(n41) );
  CIVX1 U235 ( .A(n152), .Z(n151) );
  CANR1X1 U236 ( .A(n161), .B(n153), .C(n154), .Z(n152) );
  CANR1XL U237 ( .A(n306), .B(n54), .C(n51), .Z(n49) );
  CANR1XL U238 ( .A(n305), .B(n62), .C(n59), .Z(n57) );
  CAN2X1 U239 ( .A(n299), .B(n165), .Z(SUM[0]) );
  CNIVX1 U240 ( .A(n308), .Z(SUM[1]) );
  COND1X1 U241 ( .A(n132), .B(n152), .C(n133), .Z(n131) );
  COND1X1 U242 ( .A(n55), .B(n57), .C(n56), .Z(n54) );
  CND2XL U243 ( .A(A[6]), .B(B[6]), .Z(n140) );
  CANR1XL U244 ( .A(n143), .B(n134), .C(n135), .Z(n133) );
  COND1XL U245 ( .A(n165), .B(n162), .C(n163), .Z(n161) );
  CND2XL U246 ( .A(n193), .B(n163), .Z(n28) );
  CNR2X1 U247 ( .A(A[12]), .B(B[12]), .Z(n105) );
  COND1X1 U248 ( .A(n47), .B(n49), .C(n48), .Z(n46) );
  CND2XL U249 ( .A(n142), .B(n134), .Z(n132) );
  CNR2XL U250 ( .A(n139), .B(n136), .Z(n134) );
  CNR2XL U251 ( .A(n105), .B(n100), .Z(n98) );
  CNR2XL U252 ( .A(n128), .B(n125), .Z(n123) );
  CND2IX1 U253 ( .B(n39), .A(n40), .Z(n3) );
  CND2IX1 U254 ( .B(n47), .A(n48), .Z(n5) );
  CND2IX1 U255 ( .B(n55), .A(n56), .Z(n7) );
  CNR2XL U256 ( .A(n93), .B(n88), .Z(n86) );
  CNR2XL U257 ( .A(n118), .B(n113), .Z(n111) );
  CND2IX1 U258 ( .B(n63), .A(n64), .Z(n9) );
  CEOXL U259 ( .A(n11), .B(n73), .Z(SUM[18]) );
  CND2XL U260 ( .A(n182), .B(n106), .Z(n17) );
  CND2XL U261 ( .A(n91), .B(n94), .Z(n15) );
  CND2XL U262 ( .A(n184), .B(n119), .Z(n19) );
  CEOXL U263 ( .A(n13), .B(n81), .Z(SUM[16]) );
  CND2XL U264 ( .A(n186), .B(n129), .Z(n21) );
  CND2XL U265 ( .A(n192), .B(n159), .Z(n27) );
  CND2XL U266 ( .A(n190), .B(n150), .Z(n25) );
  CEOXL U267 ( .A(n165), .B(n28), .Z(n308) );
  CNR2XL U268 ( .A(A[8]), .B(B[8]), .Z(n128) );
  CND2XL U269 ( .A(A[1]), .B(B[1]), .Z(n163) );
  CND2XL U270 ( .A(A[3]), .B(B[3]), .Z(n156) );
  CND2XL U271 ( .A(A[9]), .B(B[9]), .Z(n126) );
  CND2XL U272 ( .A(A[11]), .B(B[11]), .Z(n114) );
  CND2XL U273 ( .A(A[7]), .B(B[7]), .Z(n137) );
  CND2XL U274 ( .A(A[13]), .B(B[13]), .Z(n101) );
  CND2XL U275 ( .A(A[5]), .B(B[5]), .Z(n145) );
  CND2XL U276 ( .A(A[15]), .B(B[15]), .Z(n89) );
  COR2XL U277 ( .A(A[0]), .B(B[0]), .Z(n299) );
  CANR1XL U278 ( .A(n131), .B(n82), .C(n83), .Z(n81) );
  CNR2X1 U279 ( .A(n109), .B(n84), .Z(n82) );
  COND1XL U280 ( .A(n84), .B(n110), .C(n85), .Z(n83) );
  CND2X1 U281 ( .A(n98), .B(n86), .Z(n84) );
  CND2X1 U282 ( .A(n123), .B(n111), .Z(n109) );
  COND1XL U283 ( .A(n96), .B(n107), .C(n97), .Z(n95) );
  COND1XL U284 ( .A(n109), .B(n130), .C(n110), .Z(n108) );
  CANR1XL U285 ( .A(n142), .B(n151), .C(n143), .Z(n141) );
  COND1XL U286 ( .A(n121), .B(n130), .C(n122), .Z(n120) );
  CNR2X1 U287 ( .A(n158), .B(n155), .Z(n153) );
  COND1XL U288 ( .A(n159), .B(n155), .C(n156), .Z(n154) );
  COND1XL U289 ( .A(n129), .B(n125), .C(n126), .Z(n124) );
  COND1XL U290 ( .A(n106), .B(n100), .C(n101), .Z(n99) );
  CANR1XL U291 ( .A(n124), .B(n111), .C(n112), .Z(n110) );
  COND1XL U292 ( .A(n119), .B(n113), .C(n114), .Z(n112) );
  CENX1 U293 ( .A(n38), .B(n2), .Z(SUM[27]) );
  CND2X1 U294 ( .A(n303), .B(n37), .Z(n2) );
  COND1XL U295 ( .A(n150), .B(n144), .C(n145), .Z(n143) );
  CANR1XL U296 ( .A(n99), .B(n86), .C(n87), .Z(n85) );
  COND1XL U297 ( .A(n94), .B(n88), .C(n89), .Z(n87) );
  COND1XL U298 ( .A(n140), .B(n136), .C(n137), .Z(n135) );
  CNR2X1 U299 ( .A(n149), .B(n144), .Z(n142) );
  CENX1 U300 ( .A(n54), .B(n6), .Z(SUM[23]) );
  CND2X1 U301 ( .A(n306), .B(n53), .Z(n6) );
  CENX1 U302 ( .A(n62), .B(n8), .Z(SUM[21]) );
  CND2X1 U303 ( .A(n305), .B(n61), .Z(n8) );
  CENX1 U304 ( .A(n46), .B(n4), .Z(SUM[25]) );
  CND2X1 U305 ( .A(n307), .B(n45), .Z(n4) );
  CND2X1 U306 ( .A(n304), .B(n69), .Z(n10) );
  CEOX1 U307 ( .A(n14), .B(n90), .Z(SUM[15]) );
  CND2X1 U308 ( .A(n179), .B(n89), .Z(n14) );
  CANR1XL U309 ( .A(n91), .B(n95), .C(n92), .Z(n90) );
  CEOX1 U310 ( .A(n24), .B(n146), .Z(SUM[5]) );
  CND2X1 U311 ( .A(n189), .B(n145), .Z(n24) );
  CANR1XL U312 ( .A(n190), .B(n151), .C(n148), .Z(n146) );
  CENX1 U313 ( .A(n138), .B(n22), .Z(SUM[7]) );
  CND2X1 U314 ( .A(n187), .B(n137), .Z(n22) );
  COND1XL U315 ( .A(n139), .B(n141), .C(n140), .Z(n138) );
  CND2X1 U316 ( .A(n302), .B(n77), .Z(n12) );
  CENX1 U317 ( .A(n95), .B(n15), .Z(SUM[14]) );
  CENX1 U318 ( .A(n120), .B(n19), .Z(SUM[10]) );
  CENX1 U319 ( .A(n127), .B(n20), .Z(SUM[9]) );
  CND2X1 U320 ( .A(n185), .B(n126), .Z(n20) );
  COND1XL U321 ( .A(n128), .B(n130), .C(n129), .Z(n127) );
  CENX1 U322 ( .A(n151), .B(n25), .Z(SUM[4]) );
  CENX1 U323 ( .A(n157), .B(n26), .Z(SUM[3]) );
  CND2X1 U324 ( .A(n191), .B(n156), .Z(n26) );
  COND1XL U325 ( .A(n158), .B(n160), .C(n159), .Z(n157) );
  CND2X1 U326 ( .A(n176), .B(n72), .Z(n11) );
  CND2X1 U327 ( .A(n178), .B(n80), .Z(n13) );
  CEOX1 U328 ( .A(n16), .B(n102), .Z(SUM[13]) );
  CND2X1 U329 ( .A(n181), .B(n101), .Z(n16) );
  CANR1XL U330 ( .A(n182), .B(n108), .C(n104), .Z(n102) );
  CEOX1 U331 ( .A(n17), .B(n107), .Z(SUM[12]) );
  CEOX1 U332 ( .A(n18), .B(n115), .Z(SUM[11]) );
  CND2X1 U333 ( .A(n183), .B(n114), .Z(n18) );
  CANR1XL U334 ( .A(n184), .B(n120), .C(n117), .Z(n115) );
  CEOX1 U335 ( .A(n21), .B(n130), .Z(SUM[8]) );
  CEOX1 U336 ( .A(n23), .B(n141), .Z(SUM[6]) );
  CND2X1 U337 ( .A(n188), .B(n140), .Z(n23) );
  CEOX1 U338 ( .A(n27), .B(n160), .Z(SUM[2]) );
  CNR2X1 U339 ( .A(A[15]), .B(B[15]), .Z(n88) );
  CNR2X1 U340 ( .A(A[13]), .B(B[13]), .Z(n100) );
  CNR2X1 U341 ( .A(A[11]), .B(B[11]), .Z(n113) );
  CNR2X1 U342 ( .A(A[9]), .B(B[9]), .Z(n125) );
  CNR2X1 U343 ( .A(A[7]), .B(B[7]), .Z(n136) );
  CNR2X1 U344 ( .A(A[5]), .B(B[5]), .Z(n144) );
  CNR2X1 U345 ( .A(A[3]), .B(B[3]), .Z(n155) );
  CNR2X1 U346 ( .A(A[6]), .B(B[6]), .Z(n139) );
  CNR2X1 U347 ( .A(A[2]), .B(B[2]), .Z(n158) );
  CNR2X1 U348 ( .A(A[14]), .B(B[14]), .Z(n93) );
  CNR2X1 U349 ( .A(A[4]), .B(B[4]), .Z(n149) );
  CNR2X1 U350 ( .A(A[10]), .B(B[10]), .Z(n118) );
  CND2X1 U351 ( .A(A[0]), .B(B[0]), .Z(n165) );
  CNR2X1 U352 ( .A(A[16]), .B(B[16]), .Z(n79) );
  CNR2X1 U353 ( .A(A[18]), .B(B[18]), .Z(n71) );
  CNR2X1 U354 ( .A(A[1]), .B(B[1]), .Z(n162) );
  CENX1 U355 ( .A(n300), .B(n30), .Z(SUM[31]) );
  CENX1 U356 ( .A(B[31]), .B(A[31]), .Z(n300) );
  CAOR1X1 U357 ( .A(n303), .B(n38), .C(n35), .Z(n301) );
  CND2X1 U358 ( .A(A[4]), .B(B[4]), .Z(n150) );
  CND2X1 U359 ( .A(A[10]), .B(B[10]), .Z(n119) );
  CND2X1 U360 ( .A(A[14]), .B(B[14]), .Z(n94) );
  CND2X1 U361 ( .A(A[12]), .B(B[12]), .Z(n106) );
  CND2X1 U362 ( .A(A[8]), .B(B[8]), .Z(n129) );
  CND2X1 U363 ( .A(A[2]), .B(B[2]), .Z(n159) );
  CND2X1 U364 ( .A(A[17]), .B(B[17]), .Z(n77) );
  CND2X1 U365 ( .A(A[16]), .B(B[16]), .Z(n80) );
  COR2X1 U366 ( .A(A[17]), .B(B[17]), .Z(n302) );
  CNR2X1 U367 ( .A(A[24]), .B(B[24]), .Z(n47) );
  CNR2X1 U368 ( .A(A[20]), .B(B[20]), .Z(n63) );
  CNR2X1 U369 ( .A(A[26]), .B(B[26]), .Z(n39) );
  CNR2X1 U370 ( .A(A[22]), .B(B[22]), .Z(n55) );
  CND2X1 U371 ( .A(A[24]), .B(B[24]), .Z(n48) );
  CND2X1 U372 ( .A(A[19]), .B(B[19]), .Z(n69) );
  CND2X1 U373 ( .A(A[21]), .B(B[21]), .Z(n61) );
  CND2X1 U374 ( .A(A[23]), .B(B[23]), .Z(n53) );
  CND2X1 U375 ( .A(A[25]), .B(B[25]), .Z(n45) );
  CND2X1 U376 ( .A(A[27]), .B(B[27]), .Z(n37) );
  COR2X1 U377 ( .A(A[27]), .B(B[27]), .Z(n303) );
  CND2X1 U378 ( .A(A[18]), .B(B[18]), .Z(n72) );
  CND2X1 U379 ( .A(A[20]), .B(B[20]), .Z(n64) );
  CND2X1 U380 ( .A(A[26]), .B(B[26]), .Z(n40) );
  CND2X1 U381 ( .A(A[22]), .B(B[22]), .Z(n56) );
  COR2X1 U382 ( .A(A[19]), .B(B[19]), .Z(n304) );
  COR2X1 U383 ( .A(A[21]), .B(B[21]), .Z(n305) );
  COR2X1 U384 ( .A(A[23]), .B(B[23]), .Z(n306) );
  COR2X1 U385 ( .A(A[25]), .B(B[25]), .Z(n307) );
  CEOXL U386 ( .A(n9), .B(n65), .Z(SUM[20]) );
  CEOXL U387 ( .A(n7), .B(n57), .Z(SUM[22]) );
  CEOXL U388 ( .A(n5), .B(n49), .Z(SUM[24]) );
  CEOXL U389 ( .A(n3), .B(n41), .Z(SUM[26]) );
  CIVX2 U390 ( .A(n99), .Z(n97) );
  CIVX2 U391 ( .A(n98), .Z(n96) );
  CIVX2 U392 ( .A(n94), .Z(n92) );
  CIVX2 U393 ( .A(n77), .Z(n75) );
  CIVX2 U394 ( .A(n69), .Z(n67) );
  CIVX2 U395 ( .A(n61), .Z(n59) );
  CIVX2 U396 ( .A(n53), .Z(n51) );
  CIVX2 U397 ( .A(n45), .Z(n43) );
  CIVX2 U398 ( .A(n37), .Z(n35) );
  CIVX2 U399 ( .A(n162), .Z(n193) );
  CIVX2 U400 ( .A(n158), .Z(n192) );
  CIVX2 U401 ( .A(n155), .Z(n191) );
  CIVX2 U402 ( .A(n144), .Z(n189) );
  CIVX2 U403 ( .A(n139), .Z(n188) );
  CIVX2 U404 ( .A(n136), .Z(n187) );
  CIVX2 U405 ( .A(n128), .Z(n186) );
  CIVX2 U406 ( .A(n125), .Z(n185) );
  CIVX2 U407 ( .A(n113), .Z(n183) );
  CIVX2 U408 ( .A(n100), .Z(n181) );
  CIVX2 U409 ( .A(n93), .Z(n91) );
  CIVX2 U410 ( .A(n88), .Z(n179) );
  CIVX2 U411 ( .A(n79), .Z(n178) );
  CIVX2 U412 ( .A(n71), .Z(n176) );
  CIVX2 U413 ( .A(n161), .Z(n160) );
  CIVX2 U414 ( .A(n150), .Z(n148) );
  CIVX2 U415 ( .A(n149), .Z(n190) );
  CIVX2 U416 ( .A(n131), .Z(n130) );
  CIVX2 U417 ( .A(n124), .Z(n122) );
  CIVX2 U418 ( .A(n123), .Z(n121) );
  CIVX2 U419 ( .A(n119), .Z(n117) );
  CIVX2 U420 ( .A(n118), .Z(n184) );
  CIVX2 U421 ( .A(n108), .Z(n107) );
  CIVX2 U422 ( .A(n106), .Z(n104) );
  CIVX2 U423 ( .A(n105), .Z(n182) );
endmodule


module calc_DW01_add_8 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n30, n31,
         n32, n35, n37, n38, n39, n40, n41, n43, n45, n46, n47, n48, n49, n51,
         n53, n54, n55, n56, n57, n59, n61, n62, n63, n64, n65, n67, n69, n70,
         n71, n72, n73, n75, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n165, n174, n179, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n309,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308;

  CFA1X1 U3 ( .A(B[30]), .B(n31), .CI(A[30]), .CO(n30), .S(SUM[30]) );
  CFA1X1 U4 ( .A(B[29]), .B(n32), .CI(A[29]), .CO(n31), .S(SUM[29]) );
  CFA1X1 U5 ( .A(B[28]), .B(n302), .CI(A[28]), .CO(n32), .S(SUM[28]) );
  COND1X1 U227 ( .A(n71), .B(n73), .C(n72), .Z(n70) );
  COND1XL U228 ( .A(n63), .B(n65), .C(n64), .Z(n62) );
  CENXL U229 ( .A(n62), .B(n8), .Z(SUM[21]) );
  CANR1X1 U230 ( .A(n306), .B(n62), .C(n59), .Z(n57) );
  CENXL U231 ( .A(n54), .B(n6), .Z(SUM[23]) );
  CANR1X1 U232 ( .A(n307), .B(n54), .C(n51), .Z(n49) );
  COND1X1 U233 ( .A(n55), .B(n57), .C(n56), .Z(n54) );
  COND1X1 U234 ( .A(n39), .B(n299), .C(n40), .Z(n38) );
  CANR1X1 U235 ( .A(n308), .B(n46), .C(n43), .Z(n299) );
  CIVXL U236 ( .A(n161), .Z(n160) );
  CANR1XL U237 ( .A(n131), .B(n82), .C(n83), .Z(n81) );
  CAN2X1 U238 ( .A(n301), .B(n165), .Z(SUM[0]) );
  CNIVX1 U239 ( .A(n309), .Z(SUM[1]) );
  COND1X1 U240 ( .A(n106), .B(n100), .C(n101), .Z(n99) );
  CND2XL U241 ( .A(A[12]), .B(B[12]), .Z(n106) );
  CNR2XL U242 ( .A(A[12]), .B(B[12]), .Z(n105) );
  CEOXL U243 ( .A(n7), .B(n57), .Z(SUM[22]) );
  CIVXL U244 ( .A(n152), .Z(n151) );
  CANR1X1 U245 ( .A(n161), .B(n153), .C(n154), .Z(n152) );
  COND1XL U246 ( .A(n165), .B(n162), .C(n163), .Z(n161) );
  CND2XL U247 ( .A(n193), .B(n163), .Z(n28) );
  CND2X1 U248 ( .A(A[6]), .B(B[6]), .Z(n140) );
  CIVXL U249 ( .A(n98), .Z(n96) );
  COND1X1 U250 ( .A(n79), .B(n81), .C(n80), .Z(n78) );
  COND1X1 U251 ( .A(n47), .B(n49), .C(n48), .Z(n46) );
  COND1X1 U252 ( .A(n132), .B(n152), .C(n133), .Z(n131) );
  CND2XL U253 ( .A(n142), .B(n134), .Z(n132) );
  CANR1X1 U254 ( .A(n143), .B(n134), .C(n135), .Z(n133) );
  CNR2XL U255 ( .A(n128), .B(n125), .Z(n123) );
  CND2IX1 U256 ( .B(n39), .A(n40), .Z(n3) );
  CND2IX1 U257 ( .B(n47), .A(n48), .Z(n5) );
  CNR2XL U258 ( .A(n93), .B(n88), .Z(n86) );
  CNR2XL U259 ( .A(n118), .B(n113), .Z(n111) );
  CND2IX1 U260 ( .B(n55), .A(n56), .Z(n7) );
  CND2IX1 U261 ( .B(n71), .A(n72), .Z(n11) );
  CEOXL U262 ( .A(n9), .B(n65), .Z(SUM[20]) );
  CND2XL U263 ( .A(n182), .B(n106), .Z(n17) );
  CND2XL U264 ( .A(n91), .B(n94), .Z(n15) );
  CND2XL U265 ( .A(n184), .B(n119), .Z(n19) );
  CND2IXL U266 ( .B(n79), .A(n80), .Z(n13) );
  CND2XL U267 ( .A(n186), .B(n129), .Z(n21) );
  CND2XL U268 ( .A(n192), .B(n159), .Z(n27) );
  CND2XL U269 ( .A(n190), .B(n150), .Z(n25) );
  CIVXL U270 ( .A(n149), .Z(n190) );
  CEOXL U271 ( .A(n165), .B(n28), .Z(n309) );
  CNR2XL U272 ( .A(A[8]), .B(B[8]), .Z(n128) );
  CENX1 U273 ( .A(n300), .B(n30), .Z(SUM[31]) );
  CENX1 U274 ( .A(B[31]), .B(A[31]), .Z(n300) );
  CND2XL U275 ( .A(A[1]), .B(B[1]), .Z(n163) );
  CND2XL U276 ( .A(A[3]), .B(B[3]), .Z(n156) );
  CND2XL U277 ( .A(A[9]), .B(B[9]), .Z(n126) );
  CND2XL U278 ( .A(A[7]), .B(B[7]), .Z(n137) );
  CND2XL U279 ( .A(A[13]), .B(B[13]), .Z(n101) );
  CND2XL U280 ( .A(A[5]), .B(B[5]), .Z(n145) );
  CND2XL U281 ( .A(A[11]), .B(B[11]), .Z(n114) );
  CND2XL U282 ( .A(A[15]), .B(B[15]), .Z(n89) );
  CND2XL U283 ( .A(A[16]), .B(B[16]), .Z(n80) );
  COR2XL U284 ( .A(A[0]), .B(B[0]), .Z(n301) );
  CNR2X1 U285 ( .A(n109), .B(n84), .Z(n82) );
  COND1XL U286 ( .A(n84), .B(n110), .C(n85), .Z(n83) );
  CND2X1 U287 ( .A(n98), .B(n86), .Z(n84) );
  CND2X1 U288 ( .A(n123), .B(n111), .Z(n109) );
  COND1XL U289 ( .A(n96), .B(n107), .C(n97), .Z(n95) );
  COND1XL U290 ( .A(n109), .B(n130), .C(n110), .Z(n108) );
  CANR1XL U291 ( .A(n142), .B(n151), .C(n143), .Z(n141) );
  COND1XL U292 ( .A(n121), .B(n130), .C(n122), .Z(n120) );
  CANR1XL U293 ( .A(n304), .B(n70), .C(n67), .Z(n65) );
  CNR2X1 U294 ( .A(n158), .B(n155), .Z(n153) );
  COND1XL U295 ( .A(n159), .B(n155), .C(n156), .Z(n154) );
  CNR2X1 U296 ( .A(n139), .B(n136), .Z(n134) );
  COND1XL U297 ( .A(n129), .B(n125), .C(n126), .Z(n124) );
  CANR1XL U298 ( .A(n124), .B(n111), .C(n112), .Z(n110) );
  COND1XL U299 ( .A(n119), .B(n113), .C(n114), .Z(n112) );
  CANR1XL U300 ( .A(n303), .B(n78), .C(n75), .Z(n73) );
  CANR1XL U301 ( .A(n308), .B(n46), .C(n43), .Z(n41) );
  CENX1 U302 ( .A(n38), .B(n2), .Z(SUM[27]) );
  CND2X1 U303 ( .A(n305), .B(n37), .Z(n2) );
  COND1XL U304 ( .A(n150), .B(n144), .C(n145), .Z(n143) );
  CANR1XL U305 ( .A(n99), .B(n86), .C(n87), .Z(n85) );
  COND1XL U306 ( .A(n94), .B(n88), .C(n89), .Z(n87) );
  CNR2X1 U307 ( .A(n105), .B(n100), .Z(n98) );
  COND1XL U308 ( .A(n140), .B(n136), .C(n137), .Z(n135) );
  CNR2X1 U309 ( .A(n149), .B(n144), .Z(n142) );
  CND2X1 U310 ( .A(n307), .B(n53), .Z(n6) );
  CENX1 U311 ( .A(n46), .B(n4), .Z(SUM[25]) );
  CND2X1 U312 ( .A(n308), .B(n45), .Z(n4) );
  CND2X1 U313 ( .A(n306), .B(n61), .Z(n8) );
  CND2X1 U314 ( .A(n174), .B(n64), .Z(n9) );
  CEOX1 U315 ( .A(n14), .B(n90), .Z(SUM[15]) );
  CND2X1 U316 ( .A(n179), .B(n89), .Z(n14) );
  CANR1XL U317 ( .A(n91), .B(n95), .C(n92), .Z(n90) );
  CEOX1 U318 ( .A(n24), .B(n146), .Z(SUM[5]) );
  CND2X1 U319 ( .A(n189), .B(n145), .Z(n24) );
  CANR1XL U320 ( .A(n190), .B(n151), .C(n148), .Z(n146) );
  CENX1 U321 ( .A(n138), .B(n22), .Z(SUM[7]) );
  CND2X1 U322 ( .A(n187), .B(n137), .Z(n22) );
  COND1XL U323 ( .A(n139), .B(n141), .C(n140), .Z(n138) );
  CENX1 U324 ( .A(n70), .B(n10), .Z(SUM[19]) );
  CND2X1 U325 ( .A(n304), .B(n69), .Z(n10) );
  CENX1 U326 ( .A(n78), .B(n12), .Z(SUM[17]) );
  CND2X1 U327 ( .A(n303), .B(n77), .Z(n12) );
  CENX1 U328 ( .A(n95), .B(n15), .Z(SUM[14]) );
  CENX1 U329 ( .A(n120), .B(n19), .Z(SUM[10]) );
  CENX1 U330 ( .A(n127), .B(n20), .Z(SUM[9]) );
  CND2X1 U331 ( .A(n185), .B(n126), .Z(n20) );
  COND1XL U332 ( .A(n128), .B(n130), .C(n129), .Z(n127) );
  CENX1 U333 ( .A(n151), .B(n25), .Z(SUM[4]) );
  CENX1 U334 ( .A(n157), .B(n26), .Z(SUM[3]) );
  CND2X1 U335 ( .A(n191), .B(n156), .Z(n26) );
  COND1XL U336 ( .A(n158), .B(n160), .C(n159), .Z(n157) );
  CEOX1 U337 ( .A(n16), .B(n102), .Z(SUM[13]) );
  CND2X1 U338 ( .A(n181), .B(n101), .Z(n16) );
  CANR1XL U339 ( .A(n182), .B(n108), .C(n104), .Z(n102) );
  CEOX1 U340 ( .A(n17), .B(n107), .Z(SUM[12]) );
  CEOX1 U341 ( .A(n18), .B(n115), .Z(SUM[11]) );
  CND2X1 U342 ( .A(n183), .B(n114), .Z(n18) );
  CANR1XL U343 ( .A(n184), .B(n120), .C(n117), .Z(n115) );
  CEOX1 U344 ( .A(n21), .B(n130), .Z(SUM[8]) );
  CEOX1 U345 ( .A(n23), .B(n141), .Z(SUM[6]) );
  CND2X1 U346 ( .A(n188), .B(n140), .Z(n23) );
  CEOX1 U347 ( .A(n27), .B(n160), .Z(SUM[2]) );
  CNR2X1 U348 ( .A(A[5]), .B(B[5]), .Z(n144) );
  CNR2X1 U349 ( .A(A[15]), .B(B[15]), .Z(n88) );
  CNR2X1 U350 ( .A(A[13]), .B(B[13]), .Z(n100) );
  CNR2X1 U351 ( .A(A[11]), .B(B[11]), .Z(n113) );
  CNR2X1 U352 ( .A(A[9]), .B(B[9]), .Z(n125) );
  CNR2X1 U353 ( .A(A[7]), .B(B[7]), .Z(n136) );
  CNR2X1 U354 ( .A(A[3]), .B(B[3]), .Z(n155) );
  CNR2X1 U355 ( .A(A[6]), .B(B[6]), .Z(n139) );
  CNR2X1 U356 ( .A(A[2]), .B(B[2]), .Z(n158) );
  CNR2X1 U357 ( .A(A[14]), .B(B[14]), .Z(n93) );
  CNR2X1 U358 ( .A(A[10]), .B(B[10]), .Z(n118) );
  CNR2X1 U359 ( .A(A[4]), .B(B[4]), .Z(n149) );
  CND2X1 U360 ( .A(A[0]), .B(B[0]), .Z(n165) );
  CNR2X1 U361 ( .A(A[16]), .B(B[16]), .Z(n79) );
  CNR2X1 U362 ( .A(A[18]), .B(B[18]), .Z(n71) );
  CNR2X1 U363 ( .A(A[1]), .B(B[1]), .Z(n162) );
  CAOR1X1 U364 ( .A(n305), .B(n38), .C(n35), .Z(n302) );
  CND2X1 U365 ( .A(A[4]), .B(B[4]), .Z(n150) );
  CND2X1 U366 ( .A(A[10]), .B(B[10]), .Z(n119) );
  CND2X1 U367 ( .A(A[14]), .B(B[14]), .Z(n94) );
  CND2X1 U368 ( .A(A[8]), .B(B[8]), .Z(n129) );
  CND2X1 U369 ( .A(A[2]), .B(B[2]), .Z(n159) );
  CND2X1 U370 ( .A(A[17]), .B(B[17]), .Z(n77) );
  CND2X1 U371 ( .A(A[19]), .B(B[19]), .Z(n69) );
  CND2X1 U372 ( .A(A[18]), .B(B[18]), .Z(n72) );
  COR2X1 U373 ( .A(A[17]), .B(B[17]), .Z(n303) );
  COR2X1 U374 ( .A(A[19]), .B(B[19]), .Z(n304) );
  CNR2X1 U375 ( .A(A[24]), .B(B[24]), .Z(n47) );
  CNR2X1 U376 ( .A(A[20]), .B(B[20]), .Z(n63) );
  CNR2X1 U377 ( .A(A[26]), .B(B[26]), .Z(n39) );
  CNR2X1 U378 ( .A(A[22]), .B(B[22]), .Z(n55) );
  CND2X1 U379 ( .A(A[24]), .B(B[24]), .Z(n48) );
  CND2X1 U380 ( .A(A[21]), .B(B[21]), .Z(n61) );
  CND2X1 U381 ( .A(A[23]), .B(B[23]), .Z(n53) );
  CND2X1 U382 ( .A(A[25]), .B(B[25]), .Z(n45) );
  CND2X1 U383 ( .A(A[27]), .B(B[27]), .Z(n37) );
  COR2X1 U384 ( .A(A[27]), .B(B[27]), .Z(n305) );
  CND2X1 U385 ( .A(A[20]), .B(B[20]), .Z(n64) );
  CND2X1 U386 ( .A(A[26]), .B(B[26]), .Z(n40) );
  CND2X1 U387 ( .A(A[22]), .B(B[22]), .Z(n56) );
  COR2X1 U388 ( .A(A[21]), .B(B[21]), .Z(n306) );
  COR2X1 U389 ( .A(A[23]), .B(B[23]), .Z(n307) );
  COR2X1 U390 ( .A(A[25]), .B(B[25]), .Z(n308) );
  CEOXL U391 ( .A(n11), .B(n73), .Z(SUM[18]) );
  CEOXL U392 ( .A(n13), .B(n81), .Z(SUM[16]) );
  CEOXL U393 ( .A(n5), .B(n49), .Z(SUM[24]) );
  CEOXL U394 ( .A(n3), .B(n41), .Z(SUM[26]) );
  CIVX2 U395 ( .A(n99), .Z(n97) );
  CIVX2 U396 ( .A(n94), .Z(n92) );
  CIVX2 U397 ( .A(n77), .Z(n75) );
  CIVX2 U398 ( .A(n69), .Z(n67) );
  CIVX2 U399 ( .A(n61), .Z(n59) );
  CIVX2 U400 ( .A(n53), .Z(n51) );
  CIVX2 U401 ( .A(n45), .Z(n43) );
  CIVX2 U402 ( .A(n37), .Z(n35) );
  CIVX2 U403 ( .A(n162), .Z(n193) );
  CIVX2 U404 ( .A(n158), .Z(n192) );
  CIVX2 U405 ( .A(n155), .Z(n191) );
  CIVX2 U406 ( .A(n144), .Z(n189) );
  CIVX2 U407 ( .A(n139), .Z(n188) );
  CIVX2 U408 ( .A(n136), .Z(n187) );
  CIVX2 U409 ( .A(n128), .Z(n186) );
  CIVX2 U410 ( .A(n125), .Z(n185) );
  CIVX2 U411 ( .A(n113), .Z(n183) );
  CIVX2 U412 ( .A(n100), .Z(n181) );
  CIVX2 U413 ( .A(n93), .Z(n91) );
  CIVX2 U414 ( .A(n88), .Z(n179) );
  CIVX2 U415 ( .A(n63), .Z(n174) );
  CIVX2 U416 ( .A(n150), .Z(n148) );
  CIVX2 U417 ( .A(n131), .Z(n130) );
  CIVX2 U418 ( .A(n124), .Z(n122) );
  CIVX2 U419 ( .A(n123), .Z(n121) );
  CIVX2 U420 ( .A(n119), .Z(n117) );
  CIVX2 U421 ( .A(n118), .Z(n184) );
  CIVX2 U422 ( .A(n108), .Z(n107) );
  CIVX2 U423 ( .A(n106), .Z(n104) );
  CIVX2 U424 ( .A(n105), .Z(n182) );
endmodule


module calc_DW01_add_9 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n30, n31,
         n32, n35, n37, n38, n39, n40, n41, n43, n45, n46, n47, n48, n49, n51,
         n53, n54, n55, n56, n57, n59, n61, n62, n63, n64, n65, n67, n69, n70,
         n71, n72, n73, n75, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n165, n172, n174, n179, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n308,
         n299, n300, n301, n302, n303, n304, n305, n306, n307;

  CFA1X1 U3 ( .A(B[30]), .B(n31), .CI(A[30]), .CO(n30), .S(SUM[30]) );
  CFA1X1 U4 ( .A(B[29]), .B(n32), .CI(A[29]), .CO(n31), .S(SUM[29]) );
  CFA1X1 U5 ( .A(B[28]), .B(n301), .CI(A[28]), .CO(n32), .S(SUM[28]) );
  CIVX2 U227 ( .A(n193), .Z(n28) );
  CNR2X2 U228 ( .A(n165), .B(n162), .Z(n161) );
  CIVX2 U229 ( .A(A[1]), .Z(n162) );
  CANR1X2 U230 ( .A(n305), .B(n46), .C(n43), .Z(n41) );
  COND1X2 U231 ( .A(n47), .B(n49), .C(n48), .Z(n46) );
  CANR1XL U232 ( .A(n124), .B(n111), .C(n112), .Z(n110) );
  COND1X1 U233 ( .A(n39), .B(n41), .C(n40), .Z(n38) );
  CAN2X1 U234 ( .A(n299), .B(n165), .Z(SUM[0]) );
  CNIVX1 U235 ( .A(n308), .Z(SUM[1]) );
  CND2XL U236 ( .A(A[0]), .B(B[0]), .Z(n165) );
  CANR1X1 U237 ( .A(n304), .B(n54), .C(n51), .Z(n49) );
  CANR1X1 U238 ( .A(n306), .B(n62), .C(n59), .Z(n57) );
  CIVXL U239 ( .A(n124), .Z(n122) );
  CIVXL U240 ( .A(n99), .Z(n97) );
  CIVXL U241 ( .A(n152), .Z(n151) );
  CANR1X1 U242 ( .A(n161), .B(n153), .C(n154), .Z(n152) );
  CNR2XL U243 ( .A(A[12]), .B(B[12]), .Z(n105) );
  CND2X1 U244 ( .A(A[6]), .B(B[6]), .Z(n140) );
  CIVXL U245 ( .A(n98), .Z(n96) );
  COND1X1 U246 ( .A(n79), .B(n81), .C(n80), .Z(n78) );
  COND1X1 U247 ( .A(n71), .B(n73), .C(n72), .Z(n70) );
  COND1X1 U248 ( .A(n63), .B(n65), .C(n64), .Z(n62) );
  COND1X1 U249 ( .A(n55), .B(n57), .C(n56), .Z(n54) );
  COND1X1 U250 ( .A(n132), .B(n152), .C(n133), .Z(n131) );
  CND2XL U251 ( .A(n142), .B(n134), .Z(n132) );
  CANR1X1 U252 ( .A(n143), .B(n134), .C(n135), .Z(n133) );
  CNR2XL U253 ( .A(n128), .B(n125), .Z(n123) );
  CND2IX1 U254 ( .B(n47), .A(n48), .Z(n5) );
  CND2IX1 U255 ( .B(n39), .A(n40), .Z(n3) );
  CNR2XL U256 ( .A(n93), .B(n88), .Z(n86) );
  CNR2XL U257 ( .A(n118), .B(n113), .Z(n111) );
  CEOXL U258 ( .A(n7), .B(n57), .Z(SUM[22]) );
  CND2IX1 U259 ( .B(n71), .A(n72), .Z(n11) );
  CND2XL U260 ( .A(n182), .B(n106), .Z(n17) );
  CEOXL U261 ( .A(n9), .B(n65), .Z(SUM[20]) );
  CND2XL U262 ( .A(n184), .B(n119), .Z(n19) );
  CND2XL U263 ( .A(n91), .B(n94), .Z(n15) );
  CND2IXL U264 ( .B(n79), .A(n80), .Z(n13) );
  CND2XL U265 ( .A(n192), .B(n159), .Z(n27) );
  CND2XL U266 ( .A(n186), .B(n129), .Z(n21) );
  CND2XL U267 ( .A(n190), .B(n150), .Z(n25) );
  CNR2XL U268 ( .A(A[8]), .B(B[8]), .Z(n128) );
  CND2XL U269 ( .A(A[3]), .B(B[3]), .Z(n156) );
  CND2XL U270 ( .A(A[9]), .B(B[9]), .Z(n126) );
  CND2XL U271 ( .A(A[5]), .B(B[5]), .Z(n145) );
  CND2XL U272 ( .A(A[7]), .B(B[7]), .Z(n137) );
  CND2XL U273 ( .A(A[13]), .B(B[13]), .Z(n101) );
  CND2XL U274 ( .A(A[11]), .B(B[11]), .Z(n114) );
  CND2XL U275 ( .A(A[15]), .B(B[15]), .Z(n89) );
  CND2XL U276 ( .A(A[16]), .B(B[16]), .Z(n80) );
  CEOXL U277 ( .A(n165), .B(n28), .Z(n308) );
  COR2XL U278 ( .A(A[0]), .B(B[0]), .Z(n299) );
  CANR1XL U279 ( .A(n131), .B(n82), .C(n83), .Z(n81) );
  CNR2X1 U280 ( .A(n109), .B(n84), .Z(n82) );
  COND1XL U281 ( .A(n84), .B(n110), .C(n85), .Z(n83) );
  CND2X1 U282 ( .A(n98), .B(n86), .Z(n84) );
  CND2X1 U283 ( .A(n123), .B(n111), .Z(n109) );
  COND1XL U284 ( .A(n96), .B(n107), .C(n97), .Z(n95) );
  COND1XL U285 ( .A(n109), .B(n130), .C(n110), .Z(n108) );
  CANR1XL U286 ( .A(n142), .B(n151), .C(n143), .Z(n141) );
  COND1XL U287 ( .A(n121), .B(n130), .C(n122), .Z(n120) );
  CANR1XL U288 ( .A(n303), .B(n70), .C(n67), .Z(n65) );
  CANR1XL U289 ( .A(n302), .B(n78), .C(n75), .Z(n73) );
  CNR2X1 U290 ( .A(n158), .B(n155), .Z(n153) );
  COND1XL U291 ( .A(n159), .B(n155), .C(n156), .Z(n154) );
  COND1XL U292 ( .A(n129), .B(n125), .C(n126), .Z(n124) );
  COND1XL U293 ( .A(n106), .B(n100), .C(n101), .Z(n99) );
  CNR2X1 U294 ( .A(n139), .B(n136), .Z(n134) );
  COND1XL U295 ( .A(n119), .B(n113), .C(n114), .Z(n112) );
  COND1XL U296 ( .A(n150), .B(n144), .C(n145), .Z(n143) );
  CANR1XL U297 ( .A(n99), .B(n86), .C(n87), .Z(n85) );
  COND1XL U298 ( .A(n94), .B(n88), .C(n89), .Z(n87) );
  CNR2X1 U299 ( .A(n105), .B(n100), .Z(n98) );
  CENX1 U300 ( .A(n38), .B(n2), .Z(SUM[27]) );
  CND2X1 U301 ( .A(n307), .B(n37), .Z(n2) );
  COND1XL U302 ( .A(n140), .B(n136), .C(n137), .Z(n135) );
  CNR2X1 U303 ( .A(n149), .B(n144), .Z(n142) );
  CENX1 U304 ( .A(n46), .B(n4), .Z(SUM[25]) );
  CND2X1 U305 ( .A(n305), .B(n45), .Z(n4) );
  CENX1 U306 ( .A(n62), .B(n8), .Z(SUM[21]) );
  CND2X1 U307 ( .A(n306), .B(n61), .Z(n8) );
  CENX1 U308 ( .A(n54), .B(n6), .Z(SUM[23]) );
  CND2X1 U309 ( .A(n304), .B(n53), .Z(n6) );
  CEOX1 U310 ( .A(n14), .B(n90), .Z(SUM[15]) );
  CND2X1 U311 ( .A(n179), .B(n89), .Z(n14) );
  CANR1XL U312 ( .A(n91), .B(n95), .C(n92), .Z(n90) );
  CND2X1 U313 ( .A(n174), .B(n64), .Z(n9) );
  CND2X1 U314 ( .A(n172), .B(n56), .Z(n7) );
  CEOX1 U315 ( .A(n24), .B(n146), .Z(SUM[5]) );
  CND2X1 U316 ( .A(n189), .B(n145), .Z(n24) );
  CANR1XL U317 ( .A(n190), .B(n151), .C(n148), .Z(n146) );
  CENX1 U318 ( .A(n138), .B(n22), .Z(SUM[7]) );
  CND2X1 U319 ( .A(n187), .B(n137), .Z(n22) );
  COND1XL U320 ( .A(n139), .B(n141), .C(n140), .Z(n138) );
  CENX1 U321 ( .A(n157), .B(n26), .Z(SUM[3]) );
  CND2X1 U322 ( .A(n191), .B(n156), .Z(n26) );
  COND1XL U323 ( .A(n158), .B(n160), .C(n159), .Z(n157) );
  CENX1 U324 ( .A(n151), .B(n25), .Z(SUM[4]) );
  CENX1 U325 ( .A(n127), .B(n20), .Z(SUM[9]) );
  CND2X1 U326 ( .A(n185), .B(n126), .Z(n20) );
  COND1XL U327 ( .A(n128), .B(n130), .C(n129), .Z(n127) );
  CENX1 U328 ( .A(n120), .B(n19), .Z(SUM[10]) );
  CENX1 U329 ( .A(n95), .B(n15), .Z(SUM[14]) );
  CENX1 U330 ( .A(n78), .B(n12), .Z(SUM[17]) );
  CND2X1 U331 ( .A(n302), .B(n77), .Z(n12) );
  CENX1 U332 ( .A(n70), .B(n10), .Z(SUM[19]) );
  CND2X1 U333 ( .A(n303), .B(n69), .Z(n10) );
  CEOX1 U334 ( .A(n27), .B(n160), .Z(SUM[2]) );
  CEOX1 U335 ( .A(n23), .B(n141), .Z(SUM[6]) );
  CND2X1 U336 ( .A(n188), .B(n140), .Z(n23) );
  CEOX1 U337 ( .A(n21), .B(n130), .Z(SUM[8]) );
  CEOX1 U338 ( .A(n18), .B(n115), .Z(SUM[11]) );
  CND2X1 U339 ( .A(n183), .B(n114), .Z(n18) );
  CANR1XL U340 ( .A(n184), .B(n120), .C(n117), .Z(n115) );
  CEOX1 U341 ( .A(n17), .B(n107), .Z(SUM[12]) );
  CEOX1 U342 ( .A(n16), .B(n102), .Z(SUM[13]) );
  CND2X1 U343 ( .A(n181), .B(n101), .Z(n16) );
  CANR1XL U344 ( .A(n182), .B(n108), .C(n104), .Z(n102) );
  CNR2X1 U345 ( .A(A[5]), .B(B[5]), .Z(n144) );
  CNR2X1 U346 ( .A(A[7]), .B(B[7]), .Z(n136) );
  CNR2X1 U347 ( .A(A[9]), .B(B[9]), .Z(n125) );
  CNR2X1 U348 ( .A(A[11]), .B(B[11]), .Z(n113) );
  CNR2X1 U349 ( .A(A[13]), .B(B[13]), .Z(n100) );
  CNR2X1 U350 ( .A(A[15]), .B(B[15]), .Z(n88) );
  CNR2X1 U351 ( .A(A[3]), .B(B[3]), .Z(n155) );
  CNR2X1 U352 ( .A(A[2]), .B(B[2]), .Z(n158) );
  CNR2X1 U353 ( .A(A[6]), .B(B[6]), .Z(n139) );
  CNR2X1 U354 ( .A(A[4]), .B(B[4]), .Z(n149) );
  CNR2X1 U355 ( .A(A[14]), .B(B[14]), .Z(n93) );
  CNR2X1 U356 ( .A(A[10]), .B(B[10]), .Z(n118) );
  CNR2X1 U357 ( .A(A[16]), .B(B[16]), .Z(n79) );
  CNR2X1 U358 ( .A(A[18]), .B(B[18]), .Z(n71) );
  CENX1 U359 ( .A(n300), .B(n30), .Z(SUM[31]) );
  CENX1 U360 ( .A(B[31]), .B(A[31]), .Z(n300) );
  CAOR1X1 U361 ( .A(n307), .B(n38), .C(n35), .Z(n301) );
  CND2X1 U362 ( .A(A[4]), .B(B[4]), .Z(n150) );
  CND2X1 U363 ( .A(A[10]), .B(B[10]), .Z(n119) );
  CND2X1 U364 ( .A(A[14]), .B(B[14]), .Z(n94) );
  CND2X1 U365 ( .A(A[12]), .B(B[12]), .Z(n106) );
  CND2X1 U366 ( .A(A[18]), .B(B[18]), .Z(n72) );
  CND2X1 U367 ( .A(A[2]), .B(B[2]), .Z(n159) );
  CND2X1 U368 ( .A(A[8]), .B(B[8]), .Z(n129) );
  CND2X1 U369 ( .A(A[17]), .B(B[17]), .Z(n77) );
  CND2X1 U370 ( .A(A[19]), .B(B[19]), .Z(n69) );
  COR2X1 U371 ( .A(A[17]), .B(B[17]), .Z(n302) );
  COR2X1 U372 ( .A(A[19]), .B(B[19]), .Z(n303) );
  CNR2X1 U373 ( .A(A[24]), .B(B[24]), .Z(n47) );
  CNR2X1 U374 ( .A(A[26]), .B(B[26]), .Z(n39) );
  CNR2X1 U375 ( .A(A[20]), .B(B[20]), .Z(n63) );
  CNR2X1 U376 ( .A(A[22]), .B(B[22]), .Z(n55) );
  CND2X1 U377 ( .A(A[24]), .B(B[24]), .Z(n48) );
  CND2X1 U378 ( .A(A[26]), .B(B[26]), .Z(n40) );
  CND2X1 U379 ( .A(A[21]), .B(B[21]), .Z(n61) );
  CND2X1 U380 ( .A(A[23]), .B(B[23]), .Z(n53) );
  CND2X1 U381 ( .A(A[25]), .B(B[25]), .Z(n45) );
  CND2X1 U382 ( .A(A[27]), .B(B[27]), .Z(n37) );
  COR2X1 U383 ( .A(A[23]), .B(B[23]), .Z(n304) );
  COR2X1 U384 ( .A(A[25]), .B(B[25]), .Z(n305) );
  CND2X1 U385 ( .A(A[20]), .B(B[20]), .Z(n64) );
  CND2X1 U386 ( .A(A[22]), .B(B[22]), .Z(n56) );
  COR2X1 U387 ( .A(A[21]), .B(B[21]), .Z(n306) );
  COR2X1 U388 ( .A(A[27]), .B(B[27]), .Z(n307) );
  CEOXL U389 ( .A(n5), .B(n49), .Z(SUM[24]) );
  CEOXL U390 ( .A(n11), .B(n73), .Z(SUM[18]) );
  CEOXL U391 ( .A(n13), .B(n81), .Z(SUM[16]) );
  CEOXL U392 ( .A(n3), .B(n41), .Z(SUM[26]) );
  CIVX2 U393 ( .A(n94), .Z(n92) );
  CIVX2 U394 ( .A(n77), .Z(n75) );
  CIVX2 U395 ( .A(n69), .Z(n67) );
  CIVX2 U396 ( .A(n61), .Z(n59) );
  CIVX2 U397 ( .A(n53), .Z(n51) );
  CIVX2 U398 ( .A(n45), .Z(n43) );
  CIVX2 U399 ( .A(n37), .Z(n35) );
  CIVX2 U400 ( .A(n162), .Z(n193) );
  CIVX2 U401 ( .A(n158), .Z(n192) );
  CIVX2 U402 ( .A(n155), .Z(n191) );
  CIVX2 U403 ( .A(n144), .Z(n189) );
  CIVX2 U404 ( .A(n139), .Z(n188) );
  CIVX2 U405 ( .A(n136), .Z(n187) );
  CIVX2 U406 ( .A(n128), .Z(n186) );
  CIVX2 U407 ( .A(n125), .Z(n185) );
  CIVX2 U408 ( .A(n113), .Z(n183) );
  CIVX2 U409 ( .A(n100), .Z(n181) );
  CIVX2 U410 ( .A(n93), .Z(n91) );
  CIVX2 U411 ( .A(n88), .Z(n179) );
  CIVX2 U412 ( .A(n63), .Z(n174) );
  CIVX2 U413 ( .A(n55), .Z(n172) );
  CIVX2 U414 ( .A(n161), .Z(n160) );
  CIVX2 U415 ( .A(n150), .Z(n148) );
  CIVX2 U416 ( .A(n149), .Z(n190) );
  CIVX2 U417 ( .A(n131), .Z(n130) );
  CIVX2 U418 ( .A(n123), .Z(n121) );
  CIVX2 U419 ( .A(n119), .Z(n117) );
  CIVX2 U420 ( .A(n118), .Z(n184) );
  CIVX2 U421 ( .A(n108), .Z(n107) );
  CIVX2 U422 ( .A(n106), .Z(n104) );
  CIVX2 U423 ( .A(n105), .Z(n182) );
endmodule


module calc_DW01_add_10 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n30, n31,
         n32, n35, n37, n38, n39, n40, n41, n43, n45, n46, n47, n48, n49, n51,
         n53, n54, n55, n56, n57, n59, n61, n62, n63, n64, n65, n67, n69, n70,
         n71, n72, n73, n75, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n165, n172, n174, n179, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308;

  CFA1X1 U3 ( .A(B[30]), .B(n31), .CI(A[30]), .CO(n30), .S(SUM[30]) );
  CFA1X1 U4 ( .A(B[29]), .B(n32), .CI(A[29]), .CO(n31), .S(SUM[29]) );
  CFA1X1 U5 ( .A(B[28]), .B(n302), .CI(A[28]), .CO(n32), .S(SUM[28]) );
  CANR1X1 U227 ( .A(n307), .B(n62), .C(n59), .Z(n57) );
  COND1XL U228 ( .A(n47), .B(n49), .C(n48), .Z(n46) );
  COND1XL U229 ( .A(n106), .B(n100), .C(n101), .Z(n99) );
  CANR1XL U230 ( .A(n143), .B(n134), .C(n135), .Z(n133) );
  CANR1X1 U231 ( .A(n305), .B(n54), .C(n51), .Z(n49) );
  CAN2XL U232 ( .A(n301), .B(n165), .Z(SUM[0]) );
  CEOX1 U233 ( .A(n165), .B(n28), .Z(SUM[1]) );
  CND2XL U234 ( .A(A[0]), .B(B[0]), .Z(n165) );
  CIVXL U235 ( .A(n99), .Z(n97) );
  CANR1X1 U236 ( .A(n303), .B(n78), .C(n75), .Z(n298) );
  CANR1X1 U237 ( .A(n306), .B(n46), .C(n43), .Z(n299) );
  CIVXL U238 ( .A(n152), .Z(n151) );
  CANR1X1 U239 ( .A(n161), .B(n153), .C(n154), .Z(n152) );
  CNR2XL U240 ( .A(A[12]), .B(B[12]), .Z(n105) );
  COND1XL U241 ( .A(n165), .B(n162), .C(n163), .Z(n161) );
  CND2XL U242 ( .A(n193), .B(n163), .Z(n28) );
  CND2X1 U243 ( .A(A[6]), .B(B[6]), .Z(n140) );
  CIVXL U244 ( .A(n98), .Z(n96) );
  COND1X1 U245 ( .A(n39), .B(n299), .C(n40), .Z(n38) );
  COND1X1 U246 ( .A(n79), .B(n81), .C(n80), .Z(n78) );
  COND1X1 U247 ( .A(n71), .B(n298), .C(n72), .Z(n70) );
  COND1X1 U248 ( .A(n63), .B(n65), .C(n64), .Z(n62) );
  COND1X1 U249 ( .A(n55), .B(n57), .C(n56), .Z(n54) );
  COND1X1 U250 ( .A(n132), .B(n152), .C(n133), .Z(n131) );
  CND2XL U251 ( .A(n142), .B(n134), .Z(n132) );
  CNR2XL U252 ( .A(n128), .B(n125), .Z(n123) );
  CND2IX1 U253 ( .B(n47), .A(n48), .Z(n5) );
  CND2IX1 U254 ( .B(n39), .A(n40), .Z(n3) );
  CNR2XL U255 ( .A(n93), .B(n88), .Z(n86) );
  CNR2XL U256 ( .A(n118), .B(n113), .Z(n111) );
  CEOXL U257 ( .A(n7), .B(n57), .Z(SUM[22]) );
  CND2IX1 U258 ( .B(n71), .A(n72), .Z(n11) );
  CND2XL U259 ( .A(n182), .B(n106), .Z(n17) );
  CEOXL U260 ( .A(n9), .B(n65), .Z(SUM[20]) );
  CND2XL U261 ( .A(n184), .B(n119), .Z(n19) );
  CND2XL U262 ( .A(n91), .B(n94), .Z(n15) );
  CND2IXL U263 ( .B(n79), .A(n80), .Z(n13) );
  CND2XL U264 ( .A(n192), .B(n159), .Z(n27) );
  CND2XL U265 ( .A(n186), .B(n129), .Z(n21) );
  CND2XL U266 ( .A(n190), .B(n150), .Z(n25) );
  CNR2XL U267 ( .A(A[8]), .B(B[8]), .Z(n128) );
  CENX1 U268 ( .A(n300), .B(n30), .Z(SUM[31]) );
  CENX1 U269 ( .A(B[31]), .B(A[31]), .Z(n300) );
  CND2XL U270 ( .A(A[1]), .B(B[1]), .Z(n163) );
  CND2XL U271 ( .A(A[3]), .B(B[3]), .Z(n156) );
  CND2XL U272 ( .A(A[9]), .B(B[9]), .Z(n126) );
  CND2XL U273 ( .A(A[7]), .B(B[7]), .Z(n137) );
  CND2XL U274 ( .A(A[13]), .B(B[13]), .Z(n101) );
  CND2XL U275 ( .A(A[5]), .B(B[5]), .Z(n145) );
  CND2XL U276 ( .A(A[11]), .B(B[11]), .Z(n114) );
  CND2XL U277 ( .A(A[15]), .B(B[15]), .Z(n89) );
  CND2XL U278 ( .A(A[16]), .B(B[16]), .Z(n80) );
  COR2XL U279 ( .A(A[0]), .B(B[0]), .Z(n301) );
  CANR1XL U280 ( .A(n131), .B(n82), .C(n83), .Z(n81) );
  CNR2X1 U281 ( .A(n109), .B(n84), .Z(n82) );
  COND1XL U282 ( .A(n84), .B(n110), .C(n85), .Z(n83) );
  CND2X1 U283 ( .A(n98), .B(n86), .Z(n84) );
  CND2X1 U284 ( .A(n123), .B(n111), .Z(n109) );
  COND1XL U285 ( .A(n96), .B(n107), .C(n97), .Z(n95) );
  COND1XL U286 ( .A(n109), .B(n130), .C(n110), .Z(n108) );
  CANR1XL U287 ( .A(n142), .B(n151), .C(n143), .Z(n141) );
  COND1XL U288 ( .A(n121), .B(n130), .C(n122), .Z(n120) );
  CANR1XL U289 ( .A(n304), .B(n70), .C(n67), .Z(n65) );
  CANR1XL U290 ( .A(n303), .B(n78), .C(n75), .Z(n73) );
  CNR2X1 U291 ( .A(n158), .B(n155), .Z(n153) );
  COND1XL U292 ( .A(n159), .B(n155), .C(n156), .Z(n154) );
  COND1XL U293 ( .A(n129), .B(n125), .C(n126), .Z(n124) );
  CNR2X1 U294 ( .A(n139), .B(n136), .Z(n134) );
  CANR1XL U295 ( .A(n124), .B(n111), .C(n112), .Z(n110) );
  COND1XL U296 ( .A(n119), .B(n113), .C(n114), .Z(n112) );
  CANR1XL U297 ( .A(n306), .B(n46), .C(n43), .Z(n41) );
  COND1XL U298 ( .A(n150), .B(n144), .C(n145), .Z(n143) );
  CANR1XL U299 ( .A(n99), .B(n86), .C(n87), .Z(n85) );
  COND1XL U300 ( .A(n94), .B(n88), .C(n89), .Z(n87) );
  CNR2X1 U301 ( .A(n105), .B(n100), .Z(n98) );
  CENX1 U302 ( .A(n38), .B(n2), .Z(SUM[27]) );
  CND2X1 U303 ( .A(n308), .B(n37), .Z(n2) );
  COND1XL U304 ( .A(n140), .B(n136), .C(n137), .Z(n135) );
  CNR2X1 U305 ( .A(n149), .B(n144), .Z(n142) );
  CENX1 U306 ( .A(n46), .B(n4), .Z(SUM[25]) );
  CND2X1 U307 ( .A(n306), .B(n45), .Z(n4) );
  CENX1 U308 ( .A(n62), .B(n8), .Z(SUM[21]) );
  CND2X1 U309 ( .A(n307), .B(n61), .Z(n8) );
  CENX1 U310 ( .A(n54), .B(n6), .Z(SUM[23]) );
  CND2X1 U311 ( .A(n305), .B(n53), .Z(n6) );
  CEOX1 U312 ( .A(n14), .B(n90), .Z(SUM[15]) );
  CND2X1 U313 ( .A(n179), .B(n89), .Z(n14) );
  CANR1XL U314 ( .A(n91), .B(n95), .C(n92), .Z(n90) );
  CND2X1 U315 ( .A(n174), .B(n64), .Z(n9) );
  CND2X1 U316 ( .A(n172), .B(n56), .Z(n7) );
  CEOX1 U317 ( .A(n24), .B(n146), .Z(SUM[5]) );
  CND2X1 U318 ( .A(n189), .B(n145), .Z(n24) );
  CANR1XL U319 ( .A(n190), .B(n151), .C(n148), .Z(n146) );
  CENX1 U320 ( .A(n138), .B(n22), .Z(SUM[7]) );
  CND2X1 U321 ( .A(n187), .B(n137), .Z(n22) );
  COND1XL U322 ( .A(n139), .B(n141), .C(n140), .Z(n138) );
  CENX1 U323 ( .A(n157), .B(n26), .Z(SUM[3]) );
  CND2X1 U324 ( .A(n191), .B(n156), .Z(n26) );
  COND1XL U325 ( .A(n158), .B(n160), .C(n159), .Z(n157) );
  CENX1 U326 ( .A(n151), .B(n25), .Z(SUM[4]) );
  CENX1 U327 ( .A(n127), .B(n20), .Z(SUM[9]) );
  CND2X1 U328 ( .A(n185), .B(n126), .Z(n20) );
  COND1XL U329 ( .A(n128), .B(n130), .C(n129), .Z(n127) );
  CENX1 U330 ( .A(n120), .B(n19), .Z(SUM[10]) );
  CENX1 U331 ( .A(n95), .B(n15), .Z(SUM[14]) );
  CENX1 U332 ( .A(n78), .B(n12), .Z(SUM[17]) );
  CND2X1 U333 ( .A(n303), .B(n77), .Z(n12) );
  CENX1 U334 ( .A(n70), .B(n10), .Z(SUM[19]) );
  CND2X1 U335 ( .A(n304), .B(n69), .Z(n10) );
  CEOX1 U336 ( .A(n27), .B(n160), .Z(SUM[2]) );
  CEOX1 U337 ( .A(n23), .B(n141), .Z(SUM[6]) );
  CND2X1 U338 ( .A(n188), .B(n140), .Z(n23) );
  CEOX1 U339 ( .A(n21), .B(n130), .Z(SUM[8]) );
  CEOX1 U340 ( .A(n18), .B(n115), .Z(SUM[11]) );
  CND2X1 U341 ( .A(n183), .B(n114), .Z(n18) );
  CANR1XL U342 ( .A(n184), .B(n120), .C(n117), .Z(n115) );
  CEOX1 U343 ( .A(n17), .B(n107), .Z(SUM[12]) );
  CEOX1 U344 ( .A(n16), .B(n102), .Z(SUM[13]) );
  CND2X1 U345 ( .A(n181), .B(n101), .Z(n16) );
  CANR1XL U346 ( .A(n182), .B(n108), .C(n104), .Z(n102) );
  CNR2X1 U347 ( .A(A[5]), .B(B[5]), .Z(n144) );
  CNR2X1 U348 ( .A(A[7]), .B(B[7]), .Z(n136) );
  CNR2X1 U349 ( .A(A[9]), .B(B[9]), .Z(n125) );
  CNR2X1 U350 ( .A(A[11]), .B(B[11]), .Z(n113) );
  CNR2X1 U351 ( .A(A[13]), .B(B[13]), .Z(n100) );
  CNR2X1 U352 ( .A(A[15]), .B(B[15]), .Z(n88) );
  CNR2X1 U353 ( .A(A[3]), .B(B[3]), .Z(n155) );
  CNR2X1 U354 ( .A(A[2]), .B(B[2]), .Z(n158) );
  CNR2X1 U355 ( .A(A[6]), .B(B[6]), .Z(n139) );
  CNR2X1 U356 ( .A(A[4]), .B(B[4]), .Z(n149) );
  CNR2X1 U357 ( .A(A[14]), .B(B[14]), .Z(n93) );
  CNR2X1 U358 ( .A(A[10]), .B(B[10]), .Z(n118) );
  CNR2X1 U359 ( .A(A[16]), .B(B[16]), .Z(n79) );
  CNR2X1 U360 ( .A(A[18]), .B(B[18]), .Z(n71) );
  CNR2X1 U361 ( .A(A[1]), .B(B[1]), .Z(n162) );
  CAOR1X1 U362 ( .A(n308), .B(n38), .C(n35), .Z(n302) );
  CND2X1 U363 ( .A(A[4]), .B(B[4]), .Z(n150) );
  CND2X1 U364 ( .A(A[10]), .B(B[10]), .Z(n119) );
  CND2X1 U365 ( .A(A[14]), .B(B[14]), .Z(n94) );
  CND2X1 U366 ( .A(A[12]), .B(B[12]), .Z(n106) );
  CND2X1 U367 ( .A(A[18]), .B(B[18]), .Z(n72) );
  CND2X1 U368 ( .A(A[2]), .B(B[2]), .Z(n159) );
  CND2X1 U369 ( .A(A[8]), .B(B[8]), .Z(n129) );
  CND2X1 U370 ( .A(A[17]), .B(B[17]), .Z(n77) );
  CND2X1 U371 ( .A(A[19]), .B(B[19]), .Z(n69) );
  COR2X1 U372 ( .A(A[17]), .B(B[17]), .Z(n303) );
  COR2X1 U373 ( .A(A[19]), .B(B[19]), .Z(n304) );
  CNR2X1 U374 ( .A(A[24]), .B(B[24]), .Z(n47) );
  CNR2X1 U375 ( .A(A[26]), .B(B[26]), .Z(n39) );
  CNR2X1 U376 ( .A(A[20]), .B(B[20]), .Z(n63) );
  CNR2X1 U377 ( .A(A[22]), .B(B[22]), .Z(n55) );
  CND2X1 U378 ( .A(A[24]), .B(B[24]), .Z(n48) );
  CND2X1 U379 ( .A(A[26]), .B(B[26]), .Z(n40) );
  CND2X1 U380 ( .A(A[21]), .B(B[21]), .Z(n61) );
  CND2X1 U381 ( .A(A[23]), .B(B[23]), .Z(n53) );
  CND2X1 U382 ( .A(A[25]), .B(B[25]), .Z(n45) );
  CND2X1 U383 ( .A(A[27]), .B(B[27]), .Z(n37) );
  COR2X1 U384 ( .A(A[23]), .B(B[23]), .Z(n305) );
  COR2X1 U385 ( .A(A[25]), .B(B[25]), .Z(n306) );
  CND2X1 U386 ( .A(A[20]), .B(B[20]), .Z(n64) );
  CND2X1 U387 ( .A(A[22]), .B(B[22]), .Z(n56) );
  COR2X1 U388 ( .A(A[21]), .B(B[21]), .Z(n307) );
  COR2X1 U389 ( .A(A[27]), .B(B[27]), .Z(n308) );
  CEOXL U390 ( .A(n5), .B(n49), .Z(SUM[24]) );
  CEOXL U391 ( .A(n11), .B(n73), .Z(SUM[18]) );
  CEOXL U392 ( .A(n13), .B(n81), .Z(SUM[16]) );
  CEOXL U393 ( .A(n3), .B(n41), .Z(SUM[26]) );
  CIVX2 U394 ( .A(n94), .Z(n92) );
  CIVX2 U395 ( .A(n77), .Z(n75) );
  CIVX2 U396 ( .A(n69), .Z(n67) );
  CIVX2 U397 ( .A(n61), .Z(n59) );
  CIVX2 U398 ( .A(n53), .Z(n51) );
  CIVX2 U399 ( .A(n45), .Z(n43) );
  CIVX2 U400 ( .A(n37), .Z(n35) );
  CIVX2 U401 ( .A(n162), .Z(n193) );
  CIVX2 U402 ( .A(n158), .Z(n192) );
  CIVX2 U403 ( .A(n155), .Z(n191) );
  CIVX2 U404 ( .A(n144), .Z(n189) );
  CIVX2 U405 ( .A(n139), .Z(n188) );
  CIVX2 U406 ( .A(n136), .Z(n187) );
  CIVX2 U407 ( .A(n128), .Z(n186) );
  CIVX2 U408 ( .A(n125), .Z(n185) );
  CIVX2 U409 ( .A(n113), .Z(n183) );
  CIVX2 U410 ( .A(n100), .Z(n181) );
  CIVX2 U411 ( .A(n93), .Z(n91) );
  CIVX2 U412 ( .A(n88), .Z(n179) );
  CIVX2 U413 ( .A(n63), .Z(n174) );
  CIVX2 U414 ( .A(n55), .Z(n172) );
  CIVX2 U415 ( .A(n161), .Z(n160) );
  CIVX2 U416 ( .A(n150), .Z(n148) );
  CIVX2 U417 ( .A(n149), .Z(n190) );
  CIVX2 U418 ( .A(n131), .Z(n130) );
  CIVX2 U419 ( .A(n124), .Z(n122) );
  CIVX2 U420 ( .A(n123), .Z(n121) );
  CIVX2 U421 ( .A(n119), .Z(n117) );
  CIVX2 U422 ( .A(n118), .Z(n184) );
  CIVX2 U423 ( .A(n108), .Z(n107) );
  CIVX2 U424 ( .A(n106), .Z(n104) );
  CIVX2 U425 ( .A(n105), .Z(n182) );
endmodule


module calc_DW01_add_11 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n30, n31,
         n32, n35, n37, n38, n39, n40, n41, n43, n45, n46, n47, n48, n49, n51,
         n53, n54, n55, n56, n57, n59, n61, n62, n63, n64, n65, n67, n69, n70,
         n71, n72, n73, n75, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n165, n176, n178, n179, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n308, n299, n300, n301, n302, n303, n304, n305, n306, n307;

  CFA1X1 U3 ( .A(B[30]), .B(n31), .CI(A[30]), .CO(n30), .S(SUM[30]) );
  CFA1X1 U4 ( .A(B[29]), .B(n32), .CI(A[29]), .CO(n31), .S(SUM[29]) );
  CFA1X1 U5 ( .A(B[28]), .B(n301), .CI(A[28]), .CO(n32), .S(SUM[28]) );
  COND1X1 U58 ( .A(n63), .B(n65), .C(n64), .Z(n62) );
  CANR1X1 U227 ( .A(n307), .B(n46), .C(n43), .Z(n41) );
  CIVXL U228 ( .A(n161), .Z(n160) );
  COND1X2 U229 ( .A(n71), .B(n73), .C(n72), .Z(n70) );
  CANR1X1 U230 ( .A(n302), .B(n78), .C(n75), .Z(n73) );
  COND1X2 U231 ( .A(n55), .B(n57), .C(n56), .Z(n54) );
  CANR1X1 U232 ( .A(n305), .B(n62), .C(n59), .Z(n57) );
  COND1XL U233 ( .A(n132), .B(n152), .C(n133), .Z(n131) );
  COND1XL U234 ( .A(n39), .B(n41), .C(n40), .Z(n38) );
  CAN2X1 U235 ( .A(n299), .B(n165), .Z(SUM[0]) );
  CNIVX1 U236 ( .A(n308), .Z(SUM[1]) );
  CANR1X1 U237 ( .A(n306), .B(n54), .C(n51), .Z(n49) );
  CANR1X1 U238 ( .A(n161), .B(n153), .C(n154), .Z(n152) );
  CND2XL U239 ( .A(A[6]), .B(B[6]), .Z(n140) );
  CANR1XL U240 ( .A(n143), .B(n134), .C(n135), .Z(n133) );
  COND1XL U241 ( .A(n165), .B(n162), .C(n163), .Z(n161) );
  CND2XL U242 ( .A(n193), .B(n163), .Z(n28) );
  CNR2X1 U243 ( .A(A[12]), .B(B[12]), .Z(n105) );
  COND1X1 U244 ( .A(n79), .B(n81), .C(n80), .Z(n78) );
  COND1X1 U245 ( .A(n47), .B(n49), .C(n48), .Z(n46) );
  CND2XL U246 ( .A(n142), .B(n134), .Z(n132) );
  CNR2XL U247 ( .A(n139), .B(n136), .Z(n134) );
  CANR1X1 U248 ( .A(n304), .B(n70), .C(n67), .Z(n65) );
  CNR2XL U249 ( .A(n105), .B(n100), .Z(n98) );
  CNR2XL U250 ( .A(n128), .B(n125), .Z(n123) );
  CND2IX1 U251 ( .B(n55), .A(n56), .Z(n7) );
  CND2IX1 U252 ( .B(n47), .A(n48), .Z(n5) );
  CND2IX1 U253 ( .B(n39), .A(n40), .Z(n3) );
  CNR2XL U254 ( .A(n93), .B(n88), .Z(n86) );
  CNR2XL U255 ( .A(n118), .B(n113), .Z(n111) );
  CND2IX1 U256 ( .B(n63), .A(n64), .Z(n9) );
  CND2XL U257 ( .A(n182), .B(n106), .Z(n17) );
  CEOXL U258 ( .A(n11), .B(n73), .Z(SUM[18]) );
  CND2XL U259 ( .A(n184), .B(n119), .Z(n19) );
  CND2XL U260 ( .A(n91), .B(n94), .Z(n15) );
  CND2XL U261 ( .A(n192), .B(n159), .Z(n27) );
  CND2XL U262 ( .A(n186), .B(n129), .Z(n21) );
  CEOXL U263 ( .A(n13), .B(n81), .Z(SUM[16]) );
  CND2XL U264 ( .A(n190), .B(n150), .Z(n25) );
  CEOXL U265 ( .A(n165), .B(n28), .Z(n308) );
  CNR2XL U266 ( .A(A[8]), .B(B[8]), .Z(n128) );
  CND2XL U267 ( .A(A[1]), .B(B[1]), .Z(n163) );
  CND2XL U268 ( .A(A[3]), .B(B[3]), .Z(n156) );
  CND2XL U269 ( .A(A[9]), .B(B[9]), .Z(n126) );
  CND2XL U270 ( .A(A[11]), .B(B[11]), .Z(n114) );
  CND2XL U271 ( .A(A[7]), .B(B[7]), .Z(n137) );
  CND2XL U272 ( .A(A[13]), .B(B[13]), .Z(n101) );
  CND2XL U273 ( .A(A[5]), .B(B[5]), .Z(n145) );
  CND2XL U274 ( .A(A[15]), .B(B[15]), .Z(n89) );
  COR2XL U275 ( .A(A[0]), .B(B[0]), .Z(n299) );
  CANR1XL U276 ( .A(n131), .B(n82), .C(n83), .Z(n81) );
  CNR2X1 U277 ( .A(n109), .B(n84), .Z(n82) );
  COND1XL U278 ( .A(n84), .B(n110), .C(n85), .Z(n83) );
  CND2X1 U279 ( .A(n98), .B(n86), .Z(n84) );
  CND2X1 U280 ( .A(n123), .B(n111), .Z(n109) );
  COND1XL U281 ( .A(n96), .B(n107), .C(n97), .Z(n95) );
  COND1XL U282 ( .A(n109), .B(n130), .C(n110), .Z(n108) );
  CANR1XL U283 ( .A(n142), .B(n151), .C(n143), .Z(n141) );
  COND1XL U284 ( .A(n121), .B(n130), .C(n122), .Z(n120) );
  CNR2X1 U285 ( .A(n158), .B(n155), .Z(n153) );
  COND1XL U286 ( .A(n159), .B(n155), .C(n156), .Z(n154) );
  COND1XL U287 ( .A(n129), .B(n125), .C(n126), .Z(n124) );
  COND1XL U288 ( .A(n106), .B(n100), .C(n101), .Z(n99) );
  CANR1XL U289 ( .A(n124), .B(n111), .C(n112), .Z(n110) );
  COND1XL U290 ( .A(n119), .B(n113), .C(n114), .Z(n112) );
  CENX1 U291 ( .A(n38), .B(n2), .Z(SUM[27]) );
  CND2X1 U292 ( .A(n303), .B(n37), .Z(n2) );
  COND1XL U293 ( .A(n150), .B(n144), .C(n145), .Z(n143) );
  CANR1XL U294 ( .A(n99), .B(n86), .C(n87), .Z(n85) );
  COND1XL U295 ( .A(n94), .B(n88), .C(n89), .Z(n87) );
  COND1XL U296 ( .A(n140), .B(n136), .C(n137), .Z(n135) );
  CNR2X1 U297 ( .A(n149), .B(n144), .Z(n142) );
  CENX1 U298 ( .A(n62), .B(n8), .Z(SUM[21]) );
  CND2X1 U299 ( .A(n305), .B(n61), .Z(n8) );
  CENX1 U300 ( .A(n54), .B(n6), .Z(SUM[23]) );
  CND2X1 U301 ( .A(n306), .B(n53), .Z(n6) );
  CENX1 U302 ( .A(n70), .B(n10), .Z(SUM[19]) );
  CND2X1 U303 ( .A(n304), .B(n69), .Z(n10) );
  CENX1 U304 ( .A(n46), .B(n4), .Z(SUM[25]) );
  CND2X1 U305 ( .A(n307), .B(n45), .Z(n4) );
  CEOX1 U306 ( .A(n14), .B(n90), .Z(SUM[15]) );
  CND2X1 U307 ( .A(n179), .B(n89), .Z(n14) );
  CANR1XL U308 ( .A(n91), .B(n95), .C(n92), .Z(n90) );
  CEOX1 U309 ( .A(n24), .B(n146), .Z(SUM[5]) );
  CND2X1 U310 ( .A(n189), .B(n145), .Z(n24) );
  CANR1XL U311 ( .A(n190), .B(n151), .C(n148), .Z(n146) );
  CENX1 U312 ( .A(n138), .B(n22), .Z(SUM[7]) );
  CND2X1 U313 ( .A(n187), .B(n137), .Z(n22) );
  COND1XL U314 ( .A(n139), .B(n141), .C(n140), .Z(n138) );
  CENX1 U315 ( .A(n157), .B(n26), .Z(SUM[3]) );
  CND2X1 U316 ( .A(n191), .B(n156), .Z(n26) );
  COND1XL U317 ( .A(n158), .B(n160), .C(n159), .Z(n157) );
  CENX1 U318 ( .A(n151), .B(n25), .Z(SUM[4]) );
  CENX1 U319 ( .A(n127), .B(n20), .Z(SUM[9]) );
  CND2X1 U320 ( .A(n185), .B(n126), .Z(n20) );
  COND1XL U321 ( .A(n128), .B(n130), .C(n129), .Z(n127) );
  CENX1 U322 ( .A(n120), .B(n19), .Z(SUM[10]) );
  CENX1 U323 ( .A(n95), .B(n15), .Z(SUM[14]) );
  CENX1 U324 ( .A(n78), .B(n12), .Z(SUM[17]) );
  CND2X1 U325 ( .A(n302), .B(n77), .Z(n12) );
  CEOX1 U326 ( .A(n27), .B(n160), .Z(SUM[2]) );
  CEOX1 U327 ( .A(n23), .B(n141), .Z(SUM[6]) );
  CND2X1 U328 ( .A(n188), .B(n140), .Z(n23) );
  CEOX1 U329 ( .A(n21), .B(n130), .Z(SUM[8]) );
  CEOX1 U330 ( .A(n18), .B(n115), .Z(SUM[11]) );
  CND2X1 U331 ( .A(n183), .B(n114), .Z(n18) );
  CANR1XL U332 ( .A(n184), .B(n120), .C(n117), .Z(n115) );
  CEOX1 U333 ( .A(n17), .B(n107), .Z(SUM[12]) );
  CEOX1 U334 ( .A(n16), .B(n102), .Z(SUM[13]) );
  CND2X1 U335 ( .A(n181), .B(n101), .Z(n16) );
  CANR1XL U336 ( .A(n182), .B(n108), .C(n104), .Z(n102) );
  CND2X1 U337 ( .A(n178), .B(n80), .Z(n13) );
  CND2X1 U338 ( .A(n176), .B(n72), .Z(n11) );
  CNR2X1 U339 ( .A(A[13]), .B(B[13]), .Z(n100) );
  CNR2X1 U340 ( .A(A[15]), .B(B[15]), .Z(n88) );
  CNR2X1 U341 ( .A(A[5]), .B(B[5]), .Z(n144) );
  CNR2X1 U342 ( .A(A[7]), .B(B[7]), .Z(n136) );
  CNR2X1 U343 ( .A(A[9]), .B(B[9]), .Z(n125) );
  CNR2X1 U344 ( .A(A[11]), .B(B[11]), .Z(n113) );
  CNR2X1 U345 ( .A(A[3]), .B(B[3]), .Z(n155) );
  CNR2X1 U346 ( .A(A[2]), .B(B[2]), .Z(n158) );
  CNR2X1 U347 ( .A(A[6]), .B(B[6]), .Z(n139) );
  CNR2X1 U348 ( .A(A[14]), .B(B[14]), .Z(n93) );
  CNR2X1 U349 ( .A(A[4]), .B(B[4]), .Z(n149) );
  CNR2X1 U350 ( .A(A[10]), .B(B[10]), .Z(n118) );
  CND2X1 U351 ( .A(A[0]), .B(B[0]), .Z(n165) );
  CNR2X1 U352 ( .A(A[16]), .B(B[16]), .Z(n79) );
  CNR2X1 U353 ( .A(A[18]), .B(B[18]), .Z(n71) );
  CNR2X1 U354 ( .A(A[1]), .B(B[1]), .Z(n162) );
  CENX1 U355 ( .A(n300), .B(n30), .Z(SUM[31]) );
  CENX1 U356 ( .A(B[31]), .B(A[31]), .Z(n300) );
  CAOR1X1 U357 ( .A(n303), .B(n38), .C(n35), .Z(n301) );
  CND2X1 U358 ( .A(A[4]), .B(B[4]), .Z(n150) );
  CND2X1 U359 ( .A(A[10]), .B(B[10]), .Z(n119) );
  CND2X1 U360 ( .A(A[14]), .B(B[14]), .Z(n94) );
  CND2X1 U361 ( .A(A[12]), .B(B[12]), .Z(n106) );
  CND2X1 U362 ( .A(A[2]), .B(B[2]), .Z(n159) );
  CND2X1 U363 ( .A(A[8]), .B(B[8]), .Z(n129) );
  CND2X1 U364 ( .A(A[17]), .B(B[17]), .Z(n77) );
  CND2X1 U365 ( .A(A[16]), .B(B[16]), .Z(n80) );
  COR2X1 U366 ( .A(A[17]), .B(B[17]), .Z(n302) );
  CNR2X1 U367 ( .A(A[24]), .B(B[24]), .Z(n47) );
  CNR2X1 U368 ( .A(A[20]), .B(B[20]), .Z(n63) );
  CNR2X1 U369 ( .A(A[26]), .B(B[26]), .Z(n39) );
  CNR2X1 U370 ( .A(A[22]), .B(B[22]), .Z(n55) );
  CND2X1 U371 ( .A(A[24]), .B(B[24]), .Z(n48) );
  CND2X1 U372 ( .A(A[19]), .B(B[19]), .Z(n69) );
  CND2X1 U373 ( .A(A[21]), .B(B[21]), .Z(n61) );
  CND2X1 U374 ( .A(A[23]), .B(B[23]), .Z(n53) );
  CND2X1 U375 ( .A(A[25]), .B(B[25]), .Z(n45) );
  CND2X1 U376 ( .A(A[27]), .B(B[27]), .Z(n37) );
  COR2X1 U377 ( .A(A[27]), .B(B[27]), .Z(n303) );
  CND2X1 U378 ( .A(A[18]), .B(B[18]), .Z(n72) );
  CND2X1 U379 ( .A(A[20]), .B(B[20]), .Z(n64) );
  CND2X1 U380 ( .A(A[26]), .B(B[26]), .Z(n40) );
  CND2X1 U381 ( .A(A[22]), .B(B[22]), .Z(n56) );
  COR2X1 U382 ( .A(A[19]), .B(B[19]), .Z(n304) );
  COR2X1 U383 ( .A(A[21]), .B(B[21]), .Z(n305) );
  COR2X1 U384 ( .A(A[23]), .B(B[23]), .Z(n306) );
  COR2X1 U385 ( .A(A[25]), .B(B[25]), .Z(n307) );
  CEOXL U386 ( .A(n9), .B(n65), .Z(SUM[20]) );
  CEOXL U387 ( .A(n7), .B(n57), .Z(SUM[22]) );
  CEOXL U388 ( .A(n5), .B(n49), .Z(SUM[24]) );
  CEOXL U389 ( .A(n3), .B(n41), .Z(SUM[26]) );
  CIVX2 U390 ( .A(n99), .Z(n97) );
  CIVX2 U391 ( .A(n98), .Z(n96) );
  CIVX2 U392 ( .A(n94), .Z(n92) );
  CIVX2 U393 ( .A(n77), .Z(n75) );
  CIVX2 U394 ( .A(n69), .Z(n67) );
  CIVX2 U395 ( .A(n61), .Z(n59) );
  CIVX2 U396 ( .A(n53), .Z(n51) );
  CIVX2 U397 ( .A(n45), .Z(n43) );
  CIVX2 U398 ( .A(n37), .Z(n35) );
  CIVX2 U399 ( .A(n162), .Z(n193) );
  CIVX2 U400 ( .A(n158), .Z(n192) );
  CIVX2 U401 ( .A(n155), .Z(n191) );
  CIVX2 U402 ( .A(n144), .Z(n189) );
  CIVX2 U403 ( .A(n139), .Z(n188) );
  CIVX2 U404 ( .A(n136), .Z(n187) );
  CIVX2 U405 ( .A(n128), .Z(n186) );
  CIVX2 U406 ( .A(n125), .Z(n185) );
  CIVX2 U407 ( .A(n113), .Z(n183) );
  CIVX2 U408 ( .A(n100), .Z(n181) );
  CIVX2 U409 ( .A(n93), .Z(n91) );
  CIVX2 U410 ( .A(n88), .Z(n179) );
  CIVX2 U411 ( .A(n79), .Z(n178) );
  CIVX2 U412 ( .A(n71), .Z(n176) );
  CIVX2 U413 ( .A(n152), .Z(n151) );
  CIVX2 U414 ( .A(n150), .Z(n148) );
  CIVX2 U415 ( .A(n149), .Z(n190) );
  CIVX2 U416 ( .A(n131), .Z(n130) );
  CIVX2 U417 ( .A(n124), .Z(n122) );
  CIVX2 U418 ( .A(n123), .Z(n121) );
  CIVX2 U419 ( .A(n119), .Z(n117) );
  CIVX2 U420 ( .A(n118), .Z(n184) );
  CIVX2 U421 ( .A(n108), .Z(n107) );
  CIVX2 U422 ( .A(n106), .Z(n104) );
  CIVX2 U423 ( .A(n105), .Z(n182) );
endmodule


module calc_DW_mult_uns_11 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n6, n12, n18, n21, n24, n27, n30, n33, n36, n39, n42, n44, n48, n50,
         n53, n55, n61, n63, n66, n69, n71, n74, n77, n79, n82, n85, n87, n89,
         n91, n93, n95, n97, n99, n100, n102, n104, n105, n107, n109, n110,
         n112, n113, n114, n115, n116, n120, n122, n124, n126, n128, n130,
         n132, n134, n136, n138, n140, n142, n144, n146, n148, n150, n151,
         n152, n153, n154, n155, n156, n157, n166, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n198, n199,
         n205, n207, n208, n210, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n226, n227, n228, n229, n231, n234,
         n235, n236, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n248, n249, n250, n251, n252, n253, n257, n259, n260, n261, n262,
         n263, n269, n270, n271, n272, n273, n278, n279, n280, n281, n284,
         n285, n286, n288, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n301, n303, n304, n305, n306, n308, n311, n312, n313,
         n314, n316, n318, n319, n320, n321, n322, n323, n324, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n343, n345, n346, n348, n350, n351, n352, n354,
         n356, n357, n358, n359, n360, n362, n364, n365, n366, n367, n368,
         n370, n372, n373, n374, n375, n376, n378, n380, n382, n387, n388,
         n389, n390, n391, n393, n394, n395, n397, n399, n401, n402, n403,
         n404, n408, n410, n412, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1443, n1444,
         n1445, n1446, n1447, n1448, n1450, n1452, n1453, n1454, n1455, n1456,
         n1457, n1468, n1469, n1470, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717;
  assign n12 = a[3];
  assign n21 = a[5];
  assign n30 = a[7];
  assign n39 = a[9];
  assign n48 = a[11];
  assign n55 = a[13];
  assign n63 = a[15];
  assign n71 = a[17];
  assign n79 = a[19];
  assign n87 = a[21];
  assign n93 = a[23];
  assign n99 = a[25];
  assign n104 = a[27];
  assign n109 = a[29];
  assign n113 = a[31];
  assign n116 = b[0];
  assign n120 = b[1];
  assign n122 = b[2];
  assign n124 = b[3];
  assign n126 = b[4];
  assign n128 = b[5];
  assign n130 = b[6];
  assign n132 = b[7];
  assign n134 = b[8];
  assign n136 = b[9];
  assign n138 = b[10];
  assign n140 = b[11];
  assign n142 = b[12];
  assign n144 = b[13];
  assign n146 = b[14];
  assign n148 = b[15];
  assign n150 = b[16];
  assign n151 = b[17];
  assign n152 = b[18];
  assign n153 = b[19];
  assign n154 = b[20];
  assign n155 = b[21];
  assign n156 = b[22];
  assign n157 = b[23];

  CNR2X2 U183 ( .A(n539), .B(n562), .Z(n234) );
  COND1X1 U197 ( .A(n262), .B(n245), .C(n246), .Z(n244) );
  CNR2X2 U204 ( .A(n587), .B(n608), .Z(n249) );
  CND2X2 U205 ( .A(n587), .B(n608), .Z(n250) );
  CND2X2 U217 ( .A(n609), .B(n630), .Z(n259) );
  CNR2X2 U268 ( .A(n707), .B(n722), .Z(n295) );
  COND1X1 U292 ( .A(n330), .B(n313), .C(n314), .Z(n312) );
  CANR1X1 U294 ( .A(n1624), .B(n321), .C(n316), .Z(n314) );
  COND1X1 U304 ( .A(n328), .B(n322), .C(n323), .Z(n321) );
  CNR2X2 U307 ( .A(n767), .B(n778), .Z(n322) );
  COND1X1 U321 ( .A(n337), .B(n333), .C(n334), .Z(n332) );
  CNR2X2 U324 ( .A(n791), .B(n800), .Z(n333) );
  CEO3X2 U410 ( .A(n420), .B(n438), .C(n419), .Z(n417) );
  CEO3X2 U411 ( .A(n422), .B(n421), .C(n440), .Z(n418) );
  CEO3X2 U412 ( .A(n423), .B(n444), .C(n442), .Z(n419) );
  CEO3X2 U413 ( .A(n425), .B(n424), .C(n446), .Z(n420) );
  CEO3X2 U414 ( .A(n452), .B(n450), .C(n426), .Z(n421) );
  CEO3X2 U415 ( .A(n428), .B(n448), .C(n427), .Z(n422) );
  CEO3X2 U416 ( .A(n456), .B(n429), .C(n454), .Z(n423) );
  CEO3X2 U417 ( .A(n956), .B(n998), .C(n1106), .Z(n424) );
  CEO3X2 U418 ( .A(n938), .B(n1022), .C(n1076), .Z(n425) );
  CEO3X2 U419 ( .A(n922), .B(n976), .C(n1048), .Z(n426) );
  CEO3X2 U420 ( .A(n866), .B(n896), .C(n908), .Z(n427) );
  CEO3X2 U421 ( .A(n868), .B(n878), .C(n886), .Z(n428) );
  CFA1X1 U423 ( .A(n435), .B(n433), .CI(n460), .CO(n430), .S(n431) );
  CFA1X1 U424 ( .A(n439), .B(n462), .CI(n437), .CO(n432), .S(n433) );
  CFA1X1 U425 ( .A(n441), .B(n464), .CI(n466), .CO(n434), .S(n435) );
  CFA1X1 U426 ( .A(n443), .B(n445), .CI(n468), .CO(n436), .S(n437) );
  CFA1X1 U427 ( .A(n472), .B(n470), .CI(n447), .CO(n438), .S(n439) );
  CFA1X1 U428 ( .A(n453), .B(n449), .CI(n451), .CO(n440), .S(n441) );
  CFA1X1 U429 ( .A(n478), .B(n474), .CI(n455), .CO(n442), .S(n443) );
  CFA1X1 U430 ( .A(n480), .B(n476), .CI(n457), .CO(n444), .S(n445) );
  CFA1X1 U431 ( .A(n999), .B(n482), .CI(n484), .CO(n446), .S(n447) );
  CFA1X1 U432 ( .A(n957), .B(n1107), .CI(n1023), .CO(n448), .S(n449) );
  CFA1X1 U433 ( .A(n923), .B(n1077), .CI(n977), .CO(n450), .S(n451) );
  CFA1X1 U434 ( .A(n909), .B(n1049), .CI(n939), .CO(n452), .S(n453) );
  CFA1X1 U435 ( .A(n879), .B(n897), .CI(n1610), .CO(n454), .S(n455) );
  CFA1X1 U436 ( .A(n867), .B(n869), .CI(n873), .CO(n456), .S(n457) );
  CFA1X1 U437 ( .A(n463), .B(n461), .CI(n488), .CO(n458), .S(n459) );
  CFA1X1 U438 ( .A(n467), .B(n490), .CI(n465), .CO(n460), .S(n461) );
  CFA1X1 U439 ( .A(n469), .B(n492), .CI(n494), .CO(n462), .S(n463) );
  CFA1X1 U440 ( .A(n473), .B(n471), .CI(n496), .CO(n464), .S(n465) );
  CFA1X1 U441 ( .A(n475), .B(n498), .CI(n500), .CO(n466), .S(n467) );
  CFA1X1 U442 ( .A(n481), .B(n477), .CI(n479), .CO(n468), .S(n469) );
  CFA1X1 U443 ( .A(n502), .B(n483), .CI(n504), .CO(n470), .S(n471) );
  CFA1X1 U444 ( .A(n510), .B(n506), .CI(n508), .CO(n472), .S(n473) );
  CFA1X1 U445 ( .A(n1000), .B(n485), .CI(n1108), .CO(n474), .S(n475) );
  CFA1X1 U448 ( .A(n898), .B(n958), .CI(n910), .CO(n480), .S(n481) );
  CFA1X1 U449 ( .A(n880), .B(n888), .CI(n870), .CO(n482), .S(n483) );
  CHA1X1 U450 ( .A(n874), .B(n851), .CO(n484), .S(n485) );
  CFA1X1 U452 ( .A(n495), .B(n516), .CI(n493), .CO(n488), .S(n489) );
  CFA1X1 U453 ( .A(n497), .B(n518), .CI(n520), .CO(n490), .S(n491) );
  CFA1X1 U454 ( .A(n522), .B(n499), .CI(n501), .CO(n492), .S(n493) );
  CFA1X1 U455 ( .A(n503), .B(n524), .CI(n526), .CO(n494), .S(n495) );
  CFA1X1 U456 ( .A(n509), .B(n505), .CI(n507), .CO(n496), .S(n497) );
  CFA1X1 U457 ( .A(n511), .B(n528), .CI(n530), .CO(n498), .S(n499) );
  CFA1X1 U458 ( .A(n536), .B(n532), .CI(n534), .CO(n500), .S(n501) );
  CFA1X1 U459 ( .A(n959), .B(n1109), .CI(n1562), .CO(n502), .S(n503) );
  CFA1X1 U463 ( .A(n871), .B(n881), .CI(n875), .CO(n510), .S(n511) );
  CFA1X1 U464 ( .A(n517), .B(n515), .CI(n540), .CO(n512), .S(n513) );
  CFA1X1 U465 ( .A(n544), .B(n542), .CI(n519), .CO(n514), .S(n515) );
  CFA1X1 U466 ( .A(n546), .B(n521), .CI(n523), .CO(n516), .S(n517) );
  CFA1X1 U467 ( .A(n550), .B(n525), .CI(n548), .CO(n518), .S(n519) );
  CFA1X1 U468 ( .A(n531), .B(n527), .CI(n529), .CO(n520), .S(n521) );
  CFA1X1 U469 ( .A(n552), .B(n533), .CI(n535), .CO(n522), .S(n523) );
  CFA1X1 U470 ( .A(n558), .B(n554), .CI(n556), .CO(n524), .S(n525) );
  CFA1X1 U471 ( .A(n1002), .B(n560), .CI(n537), .CO(n526), .S(n527) );
  CFA1X1 U473 ( .A(n942), .B(n1026), .CI(n1052), .CO(n530), .S(n531) );
  CFA1X1 U475 ( .A(n876), .B(n912), .CI(n890), .CO(n534), .S(n535) );
  CHA1X1 U476 ( .A(n852), .B(n882), .CO(n536), .S(n537) );
  CFA1X1 U477 ( .A(n543), .B(n541), .CI(n564), .CO(n538), .S(n539) );
  CFA1X1 U478 ( .A(n568), .B(n545), .CI(n566), .CO(n540), .S(n541) );
  CFA1X1 U479 ( .A(n570), .B(n547), .CI(n549), .CO(n542), .S(n543) );
  CFA1X1 U480 ( .A(n574), .B(n551), .CI(n572), .CO(n544), .S(n545) );
  CFA1X1 U481 ( .A(n557), .B(n553), .CI(n555), .CO(n546), .S(n547) );
  CFA1X1 U482 ( .A(n578), .B(n559), .CI(n561), .CO(n548), .S(n549) );
  CFA1X1 U483 ( .A(n582), .B(n580), .CI(n576), .CO(n550), .S(n551) );
  CFA1X1 U484 ( .A(n1003), .B(n584), .CI(n1111), .CO(n552), .S(n553) );
  CFA1X1 U485 ( .A(n943), .B(n1053), .CI(n1027), .CO(n554), .S(n555) );
  CFA1X1 U486 ( .A(n927), .B(n1573), .CI(n1081), .CO(n556), .S(n557) );
  CFA1X1 U487 ( .A(n901), .B(n961), .CI(n913), .CO(n558), .S(n559) );
  CFA1X1 U488 ( .A(n877), .B(n1578), .CI(n883), .CO(n560), .S(n561) );
  CFA1X1 U489 ( .A(n567), .B(n565), .CI(n588), .CO(n562), .S(n563) );
  CFA1X1 U490 ( .A(n592), .B(n590), .CI(n569), .CO(n564), .S(n565) );
  CFA1X1 U491 ( .A(n594), .B(n571), .CI(n573), .CO(n566), .S(n567) );
  CFA1X1 U492 ( .A(n598), .B(n575), .CI(n596), .CO(n568), .S(n569) );
  CFA1X1 U493 ( .A(n577), .B(n581), .CI(n579), .CO(n570), .S(n571) );
  CFA1X1 U494 ( .A(n602), .B(n583), .CI(n600), .CO(n572), .S(n573) );
  CFA1X1 U495 ( .A(n585), .B(n604), .CI(n606), .CO(n574), .S(n575) );
  CFA1X1 U496 ( .A(n962), .B(n1112), .CI(n1004), .CO(n576), .S(n577) );
  CFA1X1 U497 ( .A(n944), .B(n1054), .CI(n1028), .CO(n578), .S(n579) );
  CFA1X1 U499 ( .A(n1560), .B(n914), .CI(n902), .CO(n582), .S(n583) );
  CHA1X1 U500 ( .A(n853), .B(n884), .CO(n584), .S(n585) );
  CFA1X1 U501 ( .A(n591), .B(n589), .CI(n610), .CO(n586), .S(n587) );
  CFA1X1 U502 ( .A(n614), .B(n612), .CI(n593), .CO(n588), .S(n589) );
  CFA1X1 U503 ( .A(n616), .B(n595), .CI(n597), .CO(n590), .S(n591) );
  CFA1X1 U504 ( .A(n601), .B(n599), .CI(n618), .CO(n592), .S(n593) );
  CFA1X1 U505 ( .A(n605), .B(n620), .CI(n603), .CO(n594), .S(n595) );
  CFA1X1 U506 ( .A(n624), .B(n607), .CI(n622), .CO(n596), .S(n597) );
  CFA1X1 U507 ( .A(n1005), .B(n626), .CI(n628), .CO(n598), .S(n599) );
  CFA1X1 U508 ( .A(n963), .B(n1113), .CI(n1029), .CO(n600), .S(n601) );
  CFA1X1 U509 ( .A(n1570), .B(n983), .CI(n1083), .CO(n602), .S(n603) );
  CFA1X1 U510 ( .A(n915), .B(n1558), .CI(n945), .CO(n604), .S(n605) );
  CFA1X1 U512 ( .A(n613), .B(n611), .CI(n632), .CO(n608), .S(n609) );
  CFA1X1 U513 ( .A(n617), .B(n634), .CI(n615), .CO(n610), .S(n611) );
  CFA1X1 U514 ( .A(n638), .B(n636), .CI(n619), .CO(n612), .S(n613) );
  CFA1X1 U515 ( .A(n623), .B(n640), .CI(n621), .CO(n614), .S(n615) );
  CFA1X1 U516 ( .A(n644), .B(n625), .CI(n627), .CO(n616), .S(n617) );
  CFA1X1 U517 ( .A(n648), .B(n642), .CI(n646), .CO(n618), .S(n619) );
  CFA1X1 U518 ( .A(n1006), .B(n629), .CI(n1576), .CO(n620), .S(n621) );
  CFA1X1 U519 ( .A(n964), .B(n1056), .CI(n1114), .CO(n622), .S(n623) );
  CFA1X1 U520 ( .A(n1641), .B(n984), .CI(n1084), .CO(n624), .S(n625) );
  CFA1X1 U521 ( .A(n916), .B(n946), .CI(n894), .CO(n626), .S(n627) );
  CFA1X1 U524 ( .A(n639), .B(n654), .CI(n637), .CO(n632), .S(n633) );
  CFA1X1 U525 ( .A(n658), .B(n656), .CI(n641), .CO(n634), .S(n635) );
  CFA1X1 U526 ( .A(n643), .B(n660), .CI(n645), .CO(n636), .S(n637) );
  CFA1X1 U527 ( .A(n662), .B(n647), .CI(n649), .CO(n638), .S(n639) );
  CFA1X1 U528 ( .A(n668), .B(n664), .CI(n666), .CO(n640), .S(n641) );
  CFA1X1 U529 ( .A(n965), .B(n1115), .CI(n1007), .CO(n642), .S(n643) );
  CFA1X1 U530 ( .A(n947), .B(n1031), .CI(n1085), .CO(n644), .S(n645) );
  CFA1X1 U532 ( .A(n895), .B(n917), .CI(n905), .CO(n648), .S(n649) );
  CFA1X1 U533 ( .A(n655), .B(n653), .CI(n672), .CO(n650), .S(n651) );
  CFA1X1 U534 ( .A(n659), .B(n674), .CI(n657), .CO(n652), .S(n653) );
  CFA1X1 U535 ( .A(n678), .B(n676), .CI(n661), .CO(n654), .S(n655) );
  CFA1X1 U536 ( .A(n680), .B(n663), .CI(n665), .CO(n656), .S(n657) );
  CFA1X1 U537 ( .A(n684), .B(n667), .CI(n682), .CO(n658), .S(n659) );
  CFA1X1 U538 ( .A(n1008), .B(n686), .CI(n669), .CO(n660), .S(n661) );
  CFA1X1 U539 ( .A(n986), .B(n1086), .CI(n1116), .CO(n662), .S(n663) );
  CFA1X1 U540 ( .A(n948), .B(n1032), .CI(n1058), .CO(n664), .S(n665) );
  CFA1X1 U541 ( .A(n906), .B(n932), .CI(n966), .CO(n666), .S(n667) );
  CHA1X1 U542 ( .A(n855), .B(n918), .CO(n668), .S(n669) );
  CFA1X1 U543 ( .A(n675), .B(n673), .CI(n690), .CO(n670), .S(n671) );
  CFA1X1 U544 ( .A(n679), .B(n692), .CI(n677), .CO(n672), .S(n673) );
  CFA1X1 U545 ( .A(n681), .B(n694), .CI(n696), .CO(n674), .S(n675) );
  CFA1X1 U546 ( .A(n687), .B(n683), .CI(n685), .CO(n676), .S(n677) );
  CFA1X1 U547 ( .A(n702), .B(n700), .CI(n698), .CO(n678), .S(n679) );
  CFA1X1 U548 ( .A(n987), .B(n704), .CI(n1009), .CO(n680), .S(n681) );
  CFA1X1 U549 ( .A(n967), .B(n1059), .CI(n1117), .CO(n682), .S(n683) );
  CFA1X1 U550 ( .A(n949), .B(n1087), .CI(n1033), .CO(n684), .S(n685) );
  CFA1X1 U551 ( .A(n907), .B(n933), .CI(n919), .CO(n686), .S(n687) );
  CFA1X1 U552 ( .A(n693), .B(n691), .CI(n708), .CO(n688), .S(n689) );
  CFA1X1 U553 ( .A(n697), .B(n710), .CI(n695), .CO(n690), .S(n691) );
  CFA1X1 U554 ( .A(n699), .B(n712), .CI(n714), .CO(n692), .S(n693) );
  CFA1X1 U555 ( .A(n718), .B(n701), .CI(n703), .CO(n694), .S(n695) );
  CFA1X1 U556 ( .A(n705), .B(n716), .CI(n720), .CO(n696), .S(n697) );
  CFA1X1 U557 ( .A(n988), .B(n1034), .CI(n1010), .CO(n698), .S(n699) );
  CFA1X1 U558 ( .A(n968), .B(n1088), .CI(n1118), .CO(n700), .S(n701) );
  CFA1X1 U559 ( .A(n920), .B(n934), .CI(n1060), .CO(n702), .S(n703) );
  CHA1X1 U560 ( .A(n856), .B(n950), .CO(n704), .S(n705) );
  CFA1X1 U561 ( .A(n711), .B(n709), .CI(n724), .CO(n706), .S(n707) );
  CFA1X1 U562 ( .A(n715), .B(n726), .CI(n713), .CO(n708), .S(n709) );
  CFA1X1 U563 ( .A(n717), .B(n728), .CI(n730), .CO(n710), .S(n711) );
  CFA1X1 U564 ( .A(n732), .B(n719), .CI(n721), .CO(n712), .S(n713) );
  CFA1X1 U565 ( .A(n1011), .B(n734), .CI(n736), .CO(n714), .S(n715) );
  CFA1X1 U567 ( .A(n969), .B(n1089), .CI(n1061), .CO(n718), .S(n719) );
  CFA1X1 U569 ( .A(n727), .B(n725), .CI(n740), .CO(n722), .S(n723) );
  CFA1X1 U570 ( .A(n731), .B(n742), .CI(n729), .CO(n724), .S(n725) );
  CFA1X1 U571 ( .A(n735), .B(n744), .CI(n733), .CO(n726), .S(n727) );
  CFA1X1 U572 ( .A(n750), .B(n746), .CI(n748), .CO(n728), .S(n729) );
  CFA1X1 U573 ( .A(n970), .B(n737), .CI(n1120), .CO(n730), .S(n731) );
  CFA1X1 U574 ( .A(n952), .B(n1062), .CI(n1036), .CO(n732), .S(n733) );
  CFA1X1 U575 ( .A(n936), .B(n1090), .CI(n990), .CO(n734), .S(n735) );
  CHA1X1 U576 ( .A(n857), .B(n1012), .CO(n736), .S(n737) );
  CFA1X1 U577 ( .A(n743), .B(n741), .CI(n754), .CO(n738), .S(n739) );
  CFA1X1 U578 ( .A(n758), .B(n756), .CI(n745), .CO(n740), .S(n741) );
  CFA1X1 U579 ( .A(n751), .B(n747), .CI(n749), .CO(n742), .S(n743) );
  CFA1X1 U580 ( .A(n764), .B(n762), .CI(n760), .CO(n744), .S(n745) );
  CFA1X1 U581 ( .A(n1013), .B(n1121), .CI(n1037), .CO(n746), .S(n747) );
  CFA1X1 U582 ( .A(n991), .B(n1091), .CI(n1063), .CO(n748), .S(n749) );
  CFA1X1 U583 ( .A(n971), .B(n937), .CI(n953), .CO(n750), .S(n751) );
  CFA1X1 U584 ( .A(n757), .B(n755), .CI(n768), .CO(n752), .S(n753) );
  CFA1X1 U585 ( .A(n772), .B(n759), .CI(n770), .CO(n754), .S(n755) );
  CFA1X1 U586 ( .A(n774), .B(n761), .CI(n763), .CO(n756), .S(n757) );
  CFA1X1 U587 ( .A(n992), .B(n776), .CI(n765), .CO(n758), .S(n759) );
  CFA1X1 U588 ( .A(n972), .B(n1122), .CI(n1014), .CO(n760), .S(n761) );
  CFA1X1 U589 ( .A(n954), .B(n1064), .CI(n1038), .CO(n762), .S(n763) );
  CHA1X1 U590 ( .A(n858), .B(n1092), .CO(n764), .S(n765) );
  CFA1X1 U591 ( .A(n771), .B(n769), .CI(n780), .CO(n766), .S(n767) );
  CFA1X1 U592 ( .A(n775), .B(n782), .CI(n773), .CO(n768), .S(n769) );
  CFA1X1 U593 ( .A(n784), .B(n777), .CI(n786), .CO(n770), .S(n771) );
  CFA1X1 U594 ( .A(n1039), .B(n788), .CI(n1123), .CO(n772), .S(n773) );
  CFA1X1 U595 ( .A(n1015), .B(n1065), .CI(n1093), .CO(n774), .S(n775) );
  CFA1X1 U596 ( .A(n955), .B(n993), .CI(n973), .CO(n776), .S(n777) );
  CFA1X1 U597 ( .A(n783), .B(n781), .CI(n792), .CO(n778), .S(n779) );
  CFA1X1 U598 ( .A(n787), .B(n794), .CI(n785), .CO(n780), .S(n781) );
  CFA1X1 U599 ( .A(n789), .B(n796), .CI(n798), .CO(n782), .S(n783) );
  CFA1X1 U600 ( .A(n994), .B(n1040), .CI(n1016), .CO(n784), .S(n785) );
  CFA1X1 U601 ( .A(n974), .B(n1066), .CI(n1124), .CO(n786), .S(n787) );
  CHA1X1 U602 ( .A(n859), .B(n1094), .CO(n788), .S(n789) );
  CFA1X1 U603 ( .A(n802), .B(n793), .CI(n795), .CO(n790), .S(n791) );
  CFA1X1 U604 ( .A(n799), .B(n804), .CI(n797), .CO(n792), .S(n793) );
  CFA1X1 U605 ( .A(n1125), .B(n806), .CI(n808), .CO(n794), .S(n795) );
  CFA1X1 U607 ( .A(n975), .B(n1017), .CI(n995), .CO(n798), .S(n799) );
  CFA1X1 U608 ( .A(n805), .B(n803), .CI(n812), .CO(n800), .S(n801) );
  CFA1X1 U609 ( .A(n816), .B(n807), .CI(n814), .CO(n802), .S(n803) );
  CFA1X1 U610 ( .A(n1018), .B(n809), .CI(n1042), .CO(n804), .S(n805) );
  CFA1X1 U611 ( .A(n996), .B(n1068), .CI(n1126), .CO(n806), .S(n807) );
  CHA1X1 U612 ( .A(n860), .B(n1096), .CO(n808), .S(n809) );
  CFA1X1 U613 ( .A(n815), .B(n813), .CI(n820), .CO(n810), .S(n811) );
  CFA1X1 U614 ( .A(n824), .B(n817), .CI(n822), .CO(n812), .S(n813) );
  CFA1X1 U615 ( .A(n1127), .B(n1097), .CI(n1069), .CO(n814), .S(n815) );
  CFA1X1 U616 ( .A(n997), .B(n1043), .CI(n1019), .CO(n816), .S(n817) );
  CFA1X1 U617 ( .A(n828), .B(n821), .CI(n823), .CO(n818), .S(n819) );
  CFA1X1 U618 ( .A(n1044), .B(n830), .CI(n825), .CO(n820), .S(n821) );
  CFA1X1 U619 ( .A(n1020), .B(n1070), .CI(n1128), .CO(n822), .S(n823) );
  CHA1X1 U620 ( .A(n861), .B(n1098), .CO(n824), .S(n825) );
  CFA1X1 U621 ( .A(n834), .B(n829), .CI(n831), .CO(n826), .S(n827) );
  CFA1X1 U622 ( .A(n1099), .B(n836), .CI(n1071), .CO(n828), .S(n829) );
  CFA1X1 U623 ( .A(n1021), .B(n1129), .CI(n1045), .CO(n830), .S(n831) );
  CFA1X1 U624 ( .A(n837), .B(n835), .CI(n840), .CO(n832), .S(n833) );
  CFA1X1 U625 ( .A(n1046), .B(n1072), .CI(n1130), .CO(n834), .S(n835) );
  CHA1X1 U626 ( .A(n862), .B(n1100), .CO(n836), .S(n837) );
  CFA1X1 U627 ( .A(n1073), .B(n841), .CI(n844), .CO(n838), .S(n839) );
  CFA1X1 U628 ( .A(n1566), .B(n1101), .CI(n1131), .CO(n840), .S(n841) );
  CFA1X1 U629 ( .A(n1102), .B(n845), .CI(n1074), .CO(n842), .S(n843) );
  CHA1X1 U630 ( .A(n1132), .B(n863), .CO(n844), .S(n845) );
  CFA1X1 U631 ( .A(n1565), .B(n1103), .CI(n1133), .CO(n846), .S(n847) );
  CHA1X1 U632 ( .A(n1134), .B(n1104), .CO(n848), .S(n849) );
  COND2X1 U633 ( .A(n115), .B(n1468), .C(n114), .D(n1139), .Z(n850) );
  COND2X1 U634 ( .A(n1138), .B(n115), .C(n114), .D(n1137), .Z(n866) );
  CND2IX1 U638 ( .B(n1661), .A(n113), .Z(n1139) );
  COND2X1 U639 ( .A(n112), .B(n1469), .C(n110), .D(n1144), .Z(n851) );
  COND2X1 U641 ( .A(n112), .B(n1142), .C(n110), .D(n1141), .Z(n869) );
  COND2X1 U642 ( .A(n1143), .B(n112), .C(n110), .D(n1142), .Z(n870) );
  CND2IX1 U648 ( .B(n1662), .A(n109), .Z(n1144) );
  COND2X1 U653 ( .A(n107), .B(n1149), .C(n105), .D(n1148), .Z(n875) );
  COND2X1 U654 ( .A(n1150), .B(n107), .C(n105), .D(n1149), .Z(n876) );
  CND2IX1 U662 ( .B(n1662), .A(n104), .Z(n1151) );
  COND2X1 U665 ( .A(n102), .B(n1154), .C(n1153), .D(n100), .Z(n879) );
  COND2X1 U666 ( .A(n102), .B(n1155), .C(n1154), .D(n100), .Z(n880) );
  COND2X1 U667 ( .A(n102), .B(n1156), .C(n1155), .D(n100), .Z(n881) );
  COND2X1 U668 ( .A(n102), .B(n1157), .C(n1156), .D(n100), .Z(n882) );
  COND2X1 U669 ( .A(n1158), .B(n102), .C(n1157), .D(n100), .Z(n883) );
  CND2IX1 U680 ( .B(n1662), .A(n1716), .Z(n1160) );
  COND2X1 U686 ( .A(n97), .B(n1166), .C(n1165), .D(n95), .Z(n890) );
  CND2IX1 U702 ( .B(n1662), .A(n1714), .Z(n1171) );
  COND2X1 U703 ( .A(n91), .B(n1713), .C(n1184), .D(n89), .Z(n855) );
  COND2X1 U708 ( .A(n91), .B(n1177), .C(n1176), .D(n89), .Z(n900) );
  COND2X1 U709 ( .A(n91), .B(n1178), .C(n1177), .D(n89), .Z(n901) );
  COND2X1 U710 ( .A(n91), .B(n1179), .C(n1178), .D(n89), .Z(n902) );
  COND2X1 U713 ( .A(n91), .B(n1182), .C(n1181), .D(n89), .Z(n905) );
  COND2X1 U714 ( .A(n91), .B(n1183), .C(n1182), .D(n89), .Z(n906) );
  COND2X1 U732 ( .A(n85), .B(n1188), .C(n1187), .D(n82), .Z(n910) );
  COND2X1 U734 ( .A(n85), .B(n1190), .C(n1189), .D(n82), .Z(n912) );
  COND2X1 U735 ( .A(n85), .B(n1191), .C(n1190), .D(n82), .Z(n913) );
  COND2X1 U736 ( .A(n85), .B(n1192), .C(n1191), .D(n82), .Z(n914) );
  COND2X1 U737 ( .A(n85), .B(n1193), .C(n1192), .D(n82), .Z(n915) );
  COND2X1 U738 ( .A(n85), .B(n1194), .C(n1193), .D(n82), .Z(n916) );
  COND2X1 U739 ( .A(n85), .B(n1195), .C(n1194), .D(n82), .Z(n917) );
  COND2X1 U740 ( .A(n85), .B(n1196), .C(n1195), .D(n82), .Z(n918) );
  COND2X1 U742 ( .A(n85), .B(n1198), .C(n1197), .D(n82), .Z(n920) );
  COND2X1 U765 ( .A(n77), .B(n1206), .C(n1205), .D(n74), .Z(n927) );
  COND2X1 U771 ( .A(n77), .B(n1212), .C(n1211), .D(n74), .Z(n933) );
  COND2X1 U798 ( .A(n69), .B(n1222), .C(n1221), .D(n66), .Z(n942) );
  COND2X1 U799 ( .A(n69), .B(n1223), .C(n1222), .D(n66), .Z(n943) );
  COND2X1 U800 ( .A(n69), .B(n1224), .C(n1223), .D(n66), .Z(n944) );
  COND2X1 U801 ( .A(n69), .B(n1225), .C(n1224), .D(n66), .Z(n945) );
  COND2X1 U803 ( .A(n69), .B(n1227), .C(n1226), .D(n66), .Z(n947) );
  COND2X1 U804 ( .A(n69), .B(n1228), .C(n1227), .D(n66), .Z(n948) );
  COND2X1 U805 ( .A(n69), .B(n1229), .C(n1228), .D(n66), .Z(n949) );
  COND2X1 U807 ( .A(n69), .B(n1231), .C(n1230), .D(n66), .Z(n951) );
  COND2X1 U809 ( .A(n69), .B(n1233), .C(n1232), .D(n66), .Z(n953) );
  COND2X1 U810 ( .A(n69), .B(n1234), .C(n1233), .D(n66), .Z(n954) );
  COND2X1 U832 ( .A(n61), .B(n1237), .C(n1236), .D(n1639), .Z(n956) );
  COND2X1 U833 ( .A(n61), .B(n1238), .C(n1237), .D(n1639), .Z(n957) );
  COND2X1 U834 ( .A(n61), .B(n1239), .C(n1238), .D(n1639), .Z(n958) );
  COND2X1 U835 ( .A(n61), .B(n1240), .C(n1239), .D(n1639), .Z(n959) );
  COND2X1 U836 ( .A(n61), .B(n1241), .C(n1240), .D(n1639), .Z(n960) );
  COND2X1 U838 ( .A(n61), .B(n1243), .C(n1242), .D(n1639), .Z(n962) );
  COND2X1 U839 ( .A(n61), .B(n1244), .C(n1243), .D(n1639), .Z(n963) );
  COND2X1 U840 ( .A(n61), .B(n1245), .C(n1244), .D(n1639), .Z(n964) );
  COND2X1 U841 ( .A(n61), .B(n1246), .C(n1245), .D(n1639), .Z(n965) );
  COND2X1 U844 ( .A(n61), .B(n1249), .C(n1248), .D(n1639), .Z(n968) );
  COND2X1 U845 ( .A(n61), .B(n1250), .C(n1249), .D(n1639), .Z(n969) );
  COND2X1 U846 ( .A(n61), .B(n1251), .C(n1250), .D(n1639), .Z(n970) );
  COND2X1 U847 ( .A(n61), .B(n1252), .C(n1251), .D(n1639), .Z(n971) );
  COND2X1 U848 ( .A(n61), .B(n1253), .C(n1252), .D(n1639), .Z(n972) );
  COND2X1 U849 ( .A(n61), .B(n1254), .C(n1253), .D(n1639), .Z(n973) );
  COND2X1 U850 ( .A(n61), .B(n1255), .C(n1254), .D(n1639), .Z(n974) );
  COND2X1 U883 ( .A(n53), .B(n1267), .C(n1266), .D(n50), .Z(n985) );
  COND2X1 U884 ( .A(n53), .B(n1268), .C(n1267), .D(n50), .Z(n986) );
  COND2X1 U889 ( .A(n53), .B(n1273), .C(n1272), .D(n50), .Z(n991) );
  COND2X1 U922 ( .A(n44), .B(n1283), .C(n1282), .D(n42), .Z(n1000) );
  COND2X1 U925 ( .A(n44), .B(n1286), .C(n1285), .D(n42), .Z(n1003) );
  COND2X1 U926 ( .A(n44), .B(n1287), .C(n1286), .D(n42), .Z(n1004) );
  COND2X1 U929 ( .A(n44), .B(n1290), .C(n1289), .D(n42), .Z(n1007) );
  COND2X1 U930 ( .A(n44), .B(n1291), .C(n1290), .D(n42), .Z(n1008) );
  COND2X1 U931 ( .A(n44), .B(n1292), .C(n1291), .D(n42), .Z(n1009) );
  COND2X1 U934 ( .A(n44), .B(n1295), .C(n1294), .D(n42), .Z(n1012) );
  COND2X1 U935 ( .A(n44), .B(n1296), .C(n1295), .D(n42), .Z(n1013) );
  COND2X1 U936 ( .A(n44), .B(n1297), .C(n1296), .D(n42), .Z(n1014) );
  COND2X1 U938 ( .A(n44), .B(n1299), .C(n1298), .D(n42), .Z(n1016) );
  COND2X1 U941 ( .A(n44), .B(n1302), .C(n1301), .D(n42), .Z(n1019) );
  COND2X1 U942 ( .A(n44), .B(n1303), .C(n1302), .D(n42), .Z(n1020) );
  COND2X1 U974 ( .A(n36), .B(n1310), .C(n1309), .D(n33), .Z(n1026) );
  COND2X1 U975 ( .A(n36), .B(n1311), .C(n1310), .D(n33), .Z(n1027) );
  COND2X1 U976 ( .A(n36), .B(n1312), .C(n1311), .D(n33), .Z(n1028) );
  COND2X1 U977 ( .A(n36), .B(n1313), .C(n1312), .D(n33), .Z(n1029) );
  COND2X1 U979 ( .A(n36), .B(n1315), .C(n1314), .D(n33), .Z(n1031) );
  COND2X1 U980 ( .A(n36), .B(n1316), .C(n1315), .D(n33), .Z(n1032) );
  COND2X1 U981 ( .A(n36), .B(n1317), .C(n1316), .D(n33), .Z(n1033) );
  COND2X1 U984 ( .A(n36), .B(n1320), .C(n1319), .D(n33), .Z(n1036) );
  COND2X1 U985 ( .A(n36), .B(n1321), .C(n1320), .D(n33), .Z(n1037) );
  COND2X1 U986 ( .A(n36), .B(n1322), .C(n1321), .D(n33), .Z(n1038) );
  COND2X1 U988 ( .A(n36), .B(n1324), .C(n1323), .D(n33), .Z(n1040) );
  COND2X1 U991 ( .A(n36), .B(n1327), .C(n1326), .D(n33), .Z(n1043) );
  CND2IX1 U1022 ( .B(n1661), .A(n1678), .Z(n1331) );
  COND2X1 U1033 ( .A(n27), .B(n1342), .C(n24), .D(n1341), .Z(n1057) );
  COND2X1 U1034 ( .A(n27), .B(n1343), .C(n24), .D(n1342), .Z(n1058) );
  COND2X1 U1036 ( .A(n27), .B(n1345), .C(n24), .D(n1344), .Z(n1060) );
  COND2X1 U1037 ( .A(n27), .B(n1346), .C(n24), .D(n1345), .Z(n1061) );
  COND2X1 U1039 ( .A(n27), .B(n1348), .C(n24), .D(n1347), .Z(n1063) );
  CND2IX1 U1080 ( .B(n1661), .A(n1671), .Z(n1360) );
  COND2X1 U1087 ( .A(n18), .B(n1367), .C(n1569), .D(n1366), .Z(n1081) );
  COND2X1 U1088 ( .A(n18), .B(n1368), .C(n1569), .D(n1367), .Z(n1082) );
  COND2X1 U1089 ( .A(n18), .B(n1369), .C(n1569), .D(n1368), .Z(n1083) );
  COND2X1 U1092 ( .A(n18), .B(n1372), .C(n1569), .D(n1371), .Z(n1086) );
  COND2X1 U1093 ( .A(n18), .B(n1373), .C(n1569), .D(n1372), .Z(n1087) );
  COND2X1 U1094 ( .A(n18), .B(n1374), .C(n1569), .D(n1373), .Z(n1088) );
  COND2X1 U1095 ( .A(n18), .B(n1375), .C(n1569), .D(n1374), .Z(n1089) );
  COND2X1 U1097 ( .A(n18), .B(n1377), .C(n1569), .D(n1376), .Z(n1091) );
  COND2X1 U1100 ( .A(n18), .B(n1380), .C(n1569), .D(n1379), .Z(n1094) );
  COND2X1 U1101 ( .A(n18), .B(n1381), .C(n1569), .D(n1380), .Z(n1095) );
  CND2IX1 U1142 ( .B(n1661), .A(n1664), .Z(n1391) );
  CEOX2 U1259 ( .A(a[12]), .B(n1568), .Z(n1452) );
  CEOX2 U1262 ( .A(a[10]), .B(n1694), .Z(n1453) );
  CEOX2 U1265 ( .A(a[8]), .B(n1691), .Z(n1454) );
  CEOX2 U1271 ( .A(a[4]), .B(n1676), .Z(n1456) );
  CEOX2 U1274 ( .A(a[2]), .B(n1667), .Z(n1457) );
  COND2X1 U1151 ( .A(1'b1), .B(n1400), .C(n1564), .D(n1399), .Z(n1113) );
  COND2X1 U1150 ( .A(1'b1), .B(n1399), .C(n1564), .D(n1398), .Z(n1112) );
  COND2X1 U1149 ( .A(1'b1), .B(n1398), .C(n1564), .D(n1397), .Z(n1111) );
  CNR2X2 U1281 ( .A(n1564), .B(n1392), .Z(n1106) );
  CNR2X2 U1282 ( .A(n1564), .B(n1393), .Z(n1107) );
  CNR2X2 U1283 ( .A(n1564), .B(n1394), .Z(n1108) );
  CNR2X2 U1284 ( .A(n1564), .B(n1395), .Z(n1109) );
  CNR2X2 U1285 ( .A(n1564), .B(n1396), .Z(n1110) );
  CNR2X2 U1286 ( .A(n1564), .B(n1400), .Z(n1114) );
  CNR2X2 U1287 ( .A(n1564), .B(n1413), .Z(n1127) );
  CNR2X2 U1288 ( .A(n1564), .B(n1414), .Z(n1128) );
  CNR2X2 U1289 ( .A(n1564), .B(n1415), .Z(n1129) );
  CNR2X2 U1290 ( .A(n1564), .B(n1416), .Z(n1130) );
  CNR2X2 U1291 ( .A(n1564), .B(n1417), .Z(n1131) );
  CNR2X2 U1292 ( .A(n1564), .B(n1418), .Z(n1132) );
  CNR2X2 U1293 ( .A(n1564), .B(n1419), .Z(n1133) );
  CNR2X2 U1294 ( .A(n1564), .B(n1420), .Z(n1134) );
  CNR2X2 U1295 ( .A(n1564), .B(n1421), .Z(n1135) );
  CNR2X2 U1296 ( .A(n1564), .B(n1422), .Z(n1136) );
  CNR2X2 U1297 ( .A(n1564), .B(n1412), .Z(n1126) );
  CNR2X2 U1298 ( .A(n1564), .B(n1411), .Z(n1125) );
  CNR2X2 U1299 ( .A(n1564), .B(n1410), .Z(n1124) );
  CNR2X2 U1300 ( .A(n1564), .B(n1409), .Z(n1123) );
  CNR2X2 U1301 ( .A(n1564), .B(n1408), .Z(n1122) );
  CNR2X2 U1302 ( .A(n1564), .B(n1407), .Z(n1121) );
  CNR2X2 U1303 ( .A(n1564), .B(n1406), .Z(n1120) );
  CNR2X2 U1304 ( .A(n1564), .B(n1405), .Z(n1119) );
  CNR2X2 U1305 ( .A(n1564), .B(n1404), .Z(n1118) );
  CNR2X2 U1306 ( .A(n1564), .B(n1403), .Z(n1117) );
  CNR2X2 U1307 ( .A(n1564), .B(n1402), .Z(n1116) );
  CNR2X2 U1308 ( .A(n1564), .B(n1401), .Z(n1115) );
  CIVX2 U1309 ( .A(b[31]), .Z(n1392) );
  CIVX2 U1310 ( .A(n1658), .Z(n1412) );
  CIVX2 U1311 ( .A(n1655), .Z(n1415) );
  CIVX2 U1312 ( .A(n1652), .Z(n1418) );
  CIVX2 U1313 ( .A(n1651), .Z(n1420) );
  CIVX2 U1314 ( .A(n1656), .Z(n1414) );
  CIVX2 U1315 ( .A(a[2]), .Z(n1569) );
  CIVX2 U1316 ( .A(n1649), .Z(n1422) );
  CIVX2 U1317 ( .A(n1650), .Z(n1421) );
  CIVX2 U1318 ( .A(n1657), .Z(n1413) );
  CIVX2 U1319 ( .A(n1653), .Z(n1417) );
  CIVX2 U1320 ( .A(n126), .Z(n1419) );
  CIVX2 U1321 ( .A(n148), .Z(n1408) );
  CIVX2 U1322 ( .A(n146), .Z(n1409) );
  CIVX2 U1323 ( .A(n152), .Z(n1405) );
  CENXL U1324 ( .A(1'b0), .B(n150), .Z(n1407) );
  CIVX2 U1325 ( .A(n1660), .Z(n1410) );
  CIVX2 U1326 ( .A(n1659), .Z(n1411) );
  CIVX2 U1327 ( .A(n151), .Z(n1406) );
  CIVX2 U1328 ( .A(n1136), .Z(n382) );
  CIVX2 U1329 ( .A(n382), .Z(product[1]) );
  CIVX2 U1330 ( .A(n195), .Z(product[2]) );
  CIVX2 U1331 ( .A(n378), .Z(n376) );
  CIVX2 U1332 ( .A(b[30]), .Z(n1393) );
  CIVX2 U1333 ( .A(b[29]), .Z(n1394) );
  CIVX2 U1334 ( .A(b[28]), .Z(n1395) );
  CIVX2 U1335 ( .A(b[27]), .Z(n1396) );
  CIVX2 U1336 ( .A(b[26]), .Z(n1397) );
  CIVX2 U1337 ( .A(b[25]), .Z(n1398) );
  CIVX2 U1338 ( .A(b[24]), .Z(n1399) );
  CIVX2 U1339 ( .A(n157), .Z(n1400) );
  CIVX2 U1340 ( .A(n156), .Z(n1401) );
  CIVX2 U1341 ( .A(n155), .Z(n1402) );
  CIVX2 U1342 ( .A(n154), .Z(n1403) );
  CIVX2 U1343 ( .A(n1654), .Z(n1416) );
  CIVX2 U1344 ( .A(n153), .Z(n1404) );
  COND2X1 U1346 ( .A(n97), .B(n1165), .C(n1164), .D(n95), .Z(n889) );
  CENXL U1347 ( .A(n1693), .B(n1655), .Z(n1270) );
  CENX1 U1348 ( .A(n1563), .B(n1655), .Z(n1207) );
  CENX1 U1349 ( .A(n1653), .B(n1716), .Z(n1153) );
  CENX1 U1350 ( .A(n1703), .B(n1656), .Z(n1206) );
  CNIVX1 U1351 ( .A(n1055), .Z(n1558) );
  COND1X2 U1352 ( .A(n240), .B(n234), .C(n235), .Z(n229) );
  CENX1 U1353 ( .A(n227), .B(n1577), .Z(product[27]) );
  CANR1X1 U1354 ( .A(n228), .B(n241), .C(n229), .Z(n227) );
  CANR1X1 U1355 ( .A(n279), .B(n243), .C(n244), .Z(n1559) );
  CANR1X1 U1356 ( .A(n279), .B(n243), .C(n244), .Z(n242) );
  CIVX3 U1357 ( .A(n1677), .Z(n1675) );
  CFA1X1 U1358 ( .A(n925), .B(n1051), .CI(n979), .CO(n506), .S(n507) );
  COND2X1 U1359 ( .A(n53), .B(n1261), .C(n1260), .D(n50), .Z(n979) );
  CAN2X1 U1360 ( .A(n1621), .B(n1620), .Z(n1619) );
  CIVX3 U1361 ( .A(n1715), .Z(n1714) );
  CNR2IXL U1362 ( .B(n1661), .A(n95), .Z(n895) );
  COND2X1 U1363 ( .A(n97), .B(n1170), .C(n1169), .D(n95), .Z(n894) );
  COND2X1 U1364 ( .A(n97), .B(n1163), .C(n1162), .D(n95), .Z(n887) );
  CNIVX1 U1365 ( .A(n892), .Z(n1560) );
  CIVX1 U1366 ( .A(n1001), .Z(n1561) );
  CIVX2 U1367 ( .A(n1561), .Z(n1562) );
  CFA1XL U1368 ( .A(n885), .B(n903), .CI(n893), .CO(n606), .S(n607) );
  CNIVX3 U1369 ( .A(n116), .Z(n1661) );
  COND2XL U1370 ( .A(n102), .B(n1153), .C(n1152), .D(n100), .Z(n878) );
  CIVX2 U1371 ( .A(a[16]), .Z(n1612) );
  CNIVX1 U1372 ( .A(n1702), .Z(n1563) );
  CIVXL U1373 ( .A(n1705), .Z(n1702) );
  CIVX4 U1374 ( .A(n1567), .Z(n1696) );
  CENX2 U1375 ( .A(n1716), .B(a[26]), .Z(n105) );
  CNIVX2 U1376 ( .A(n120), .Z(n1649) );
  CENXL U1377 ( .A(n1696), .B(n1657), .Z(n1245) );
  CENXL U1378 ( .A(n1708), .B(n1657), .Z(n1188) );
  CNIVX2 U1379 ( .A(n138), .Z(n1657) );
  CIVXL U1380 ( .A(n352), .Z(n351) );
  CENXL U1381 ( .A(n1674), .B(b[27]), .Z(n1332) );
  CENXL U1382 ( .A(n1674), .B(n1650), .Z(n1357) );
  CENXL U1383 ( .A(n1674), .B(n1651), .Z(n1356) );
  CENXL U1384 ( .A(n1674), .B(n1649), .Z(n1358) );
  CNIVX2 U1385 ( .A(n6), .Z(n1564) );
  COND2XL U1386 ( .A(n44), .B(n1281), .C(n1280), .D(n42), .Z(n998) );
  COND2XL U1387 ( .A(n44), .B(n1282), .C(n1281), .D(n42), .Z(n999) );
  COND2XL U1388 ( .A(n44), .B(n1294), .C(n1293), .D(n42), .Z(n1011) );
  COND2XL U1389 ( .A(n44), .B(n1301), .C(n1300), .D(n42), .Z(n1018) );
  COND2XL U1390 ( .A(n44), .B(n1285), .C(n1284), .D(n42), .Z(n1002) );
  COND2XL U1391 ( .A(n44), .B(n1293), .C(n1292), .D(n42), .Z(n1010) );
  COND2XL U1392 ( .A(n44), .B(n1289), .C(n1288), .D(n42), .Z(n1006) );
  COND2XL U1393 ( .A(n44), .B(n1300), .C(n1299), .D(n42), .Z(n1017) );
  COND2XL U1394 ( .A(n44), .B(n1288), .C(n1287), .D(n42), .Z(n1005) );
  COND2XL U1395 ( .A(n44), .B(n1284), .C(n1283), .D(n42), .Z(n1001) );
  COND2XL U1396 ( .A(n44), .B(n1298), .C(n1297), .D(n42), .Z(n1015) );
  CNIVX1 U1397 ( .A(n1075), .Z(n1565) );
  CNIVX2 U1398 ( .A(n1047), .Z(n1566) );
  CENXL U1399 ( .A(n1673), .B(n126), .Z(n1355) );
  CENXL U1400 ( .A(n1687), .B(n126), .Z(n1299) );
  CENXL U1401 ( .A(n1693), .B(n126), .Z(n1274) );
  CENXL U1402 ( .A(n1680), .B(n126), .Z(n1326) );
  CENXL U1403 ( .A(n1711), .B(n126), .Z(n1179) );
  CENXL U1404 ( .A(n1698), .B(n126), .Z(n1230) );
  CENXL U1405 ( .A(n126), .B(n104), .Z(n1146) );
  CENXL U1406 ( .A(n1696), .B(n126), .Z(n1251) );
  CENXL U1407 ( .A(n1701), .B(n126), .Z(n1211) );
  CENXL U1408 ( .A(n126), .B(n1716), .Z(n1155) );
  CENXL U1409 ( .A(n1667), .B(n126), .Z(n1386) );
  CENX1 U1410 ( .A(n1568), .B(n152), .Z(n1237) );
  CENX1 U1411 ( .A(n1563), .B(n1650), .Z(n1213) );
  CENX1 U1412 ( .A(n1696), .B(n1653), .Z(n1249) );
  CENX1 U1413 ( .A(n1696), .B(n1654), .Z(n1248) );
  CENX1 U1414 ( .A(n1671), .B(n148), .Z(n1344) );
  CENX1 U1415 ( .A(n1669), .B(n151), .Z(n1373) );
  CNR2X1 U1416 ( .A(n61), .B(n1247), .Z(n1596) );
  CENX1 U1417 ( .A(n1698), .B(n1653), .Z(n1228) );
  CENX1 U1418 ( .A(n1698), .B(n1657), .Z(n1224) );
  CENX1 U1419 ( .A(n1694), .B(n148), .Z(n1263) );
  CENX1 U1420 ( .A(n1568), .B(n1660), .Z(n1242) );
  CENX1 U1421 ( .A(n1696), .B(n1659), .Z(n1243) );
  CENX1 U1422 ( .A(n1650), .B(n1716), .Z(n1157) );
  CENX1 U1423 ( .A(n1651), .B(n1716), .Z(n1156) );
  CENX1 U1424 ( .A(n1651), .B(n104), .Z(n1147) );
  CENX1 U1425 ( .A(n1568), .B(n146), .Z(n1241) );
  CENX1 U1426 ( .A(n1698), .B(n1660), .Z(n1221) );
  CENX1 U1427 ( .A(n1697), .B(n1659), .Z(n1222) );
  CENX1 U1428 ( .A(n1568), .B(n148), .Z(n1240) );
  CENX1 U1429 ( .A(n1669), .B(n1657), .Z(n1380) );
  CENX1 U1430 ( .A(n1693), .B(n1649), .Z(n1277) );
  CENX1 U1431 ( .A(n1693), .B(n1650), .Z(n1276) );
  CENX1 U1432 ( .A(n1675), .B(n1655), .Z(n1351) );
  CENX1 U1433 ( .A(n1696), .B(n1649), .Z(n1254) );
  CENX1 U1434 ( .A(n1687), .B(n1652), .Z(n1298) );
  CENX1 U1435 ( .A(n1665), .B(n1659), .Z(n1378) );
  CENX1 U1436 ( .A(n1687), .B(n1653), .Z(n1297) );
  CENX1 U1437 ( .A(n1696), .B(n1651), .Z(n1252) );
  CENX1 U1438 ( .A(n1696), .B(n1650), .Z(n1253) );
  CENX1 U1439 ( .A(n1681), .B(n1657), .Z(n1320) );
  CENX1 U1440 ( .A(n1671), .B(n1659), .Z(n1347) );
  CENX1 U1441 ( .A(n1563), .B(n1649), .Z(n1214) );
  CENX1 U1442 ( .A(n1682), .B(n1659), .Z(n1318) );
  CENX1 U1443 ( .A(n1688), .B(n1657), .Z(n1293) );
  CENX1 U1444 ( .A(n1696), .B(n1652), .Z(n1250) );
  CENX1 U1445 ( .A(n1689), .B(n1659), .Z(n1291) );
  CENX1 U1446 ( .A(n1694), .B(n1657), .Z(n1268) );
  CENX1 U1447 ( .A(n1665), .B(n152), .Z(n1372) );
  CENX1 U1448 ( .A(n1701), .B(n1652), .Z(n1210) );
  CENX1 U1449 ( .A(n1676), .B(n151), .Z(n1342) );
  CENX1 U1450 ( .A(n1701), .B(n1653), .Z(n1209) );
  CENX1 U1451 ( .A(n1682), .B(n148), .Z(n1315) );
  CENX1 U1452 ( .A(n1697), .B(n1655), .Z(n1226) );
  CENX1 U1453 ( .A(n1683), .B(n151), .Z(n1313) );
  CENX1 U1454 ( .A(n1696), .B(n1658), .Z(n1244) );
  CENX1 U1455 ( .A(n1671), .B(n153), .Z(n1340) );
  CIVX2 U1456 ( .A(n63), .Z(n1700) );
  CENX1 U1457 ( .A(n1649), .B(n109), .Z(n1142) );
  CNIVX3 U1458 ( .A(n134), .Z(n1655) );
  CNIVX2 U1459 ( .A(n140), .Z(n1658) );
  CENX1 U1460 ( .A(n1650), .B(n109), .Z(n1141) );
  CENX1 U1461 ( .A(n1568), .B(n151), .Z(n1238) );
  CENX1 U1462 ( .A(n1678), .B(n1649), .Z(n1329) );
  CENX1 U1463 ( .A(n1687), .B(n1649), .Z(n1302) );
  CENX1 U1464 ( .A(n1680), .B(n1650), .Z(n1328) );
  CENX1 U1465 ( .A(n1673), .B(n1653), .Z(n1353) );
  CENX1 U1466 ( .A(n1687), .B(n1650), .Z(n1301) );
  CND2X2 U1467 ( .A(n1454), .B(n42), .Z(n44) );
  CIVX3 U1468 ( .A(n1635), .Z(n42) );
  CENX1 U1469 ( .A(n1685), .B(a[8]), .Z(n1635) );
  CNIVX4 U1470 ( .A(n124), .Z(n1651) );
  CENX1 U1471 ( .A(n1708), .B(n1659), .Z(n1186) );
  CENX1 U1472 ( .A(a[18]), .B(n79), .Z(n1617) );
  CENX1 U1473 ( .A(n1693), .B(n153), .Z(n1259) );
  CND2X2 U1474 ( .A(n1450), .B(n74), .Z(n77) );
  CND2X1 U1475 ( .A(n1445), .B(n105), .Z(n107) );
  CNIVX1 U1476 ( .A(n887), .Z(n1610) );
  CENX1 U1477 ( .A(n1678), .B(b[25]), .Z(n1305) );
  CENX1 U1478 ( .A(n1568), .B(n153), .Z(n1236) );
  CND2X1 U1479 ( .A(n1608), .B(n1609), .Z(n1447) );
  CENX1 U1480 ( .A(n1649), .B(n113), .Z(n1137) );
  CENX1 U1481 ( .A(n1667), .B(n1650), .Z(n1388) );
  CANR1XL U1482 ( .A(n1628), .B(n357), .C(n354), .Z(n352) );
  COND1X1 U1483 ( .A(n299), .B(n295), .C(n296), .Z(n294) );
  CNR2X1 U1484 ( .A(n631), .B(n650), .Z(n269) );
  CND2X1 U1485 ( .A(n651), .B(n670), .Z(n273) );
  CND3XL U1486 ( .A(n1645), .B(n1646), .C(n1647), .Z(n630) );
  COND1X1 U1487 ( .A(n273), .B(n269), .C(n270), .Z(n1611) );
  COND1XL U1488 ( .A(n226), .B(n218), .C(n219), .Z(n217) );
  COND1XL U1489 ( .A(n358), .B(n360), .C(n359), .Z(n357) );
  CND2X1 U1490 ( .A(n779), .B(n790), .Z(n328) );
  CIVX2 U1491 ( .A(a[0]), .Z(n6) );
  CND2X1 U1492 ( .A(n723), .B(n738), .Z(n303) );
  CND2X1 U1493 ( .A(n739), .B(n752), .Z(n306) );
  CENX1 U1494 ( .A(n241), .B(n172), .Z(product[25]) );
  CIVX2 U1495 ( .A(n1700), .Z(n1698) );
  CENX1 U1496 ( .A(n1697), .B(n1649), .Z(n1233) );
  COND2XL U1497 ( .A(n18), .B(n1379), .C(n1569), .D(n1378), .Z(n1093) );
  COND2XL U1498 ( .A(n18), .B(n1382), .C(n1569), .D(n1381), .Z(n1096) );
  CND2X1 U1499 ( .A(n1591), .B(n1592), .Z(n1085) );
  COR2X1 U1500 ( .A(n18), .B(n1371), .Z(n1591) );
  CIVX2 U1501 ( .A(n39), .Z(n1692) );
  CIVX1 U1502 ( .A(n30), .Z(n1684) );
  CIVX2 U1503 ( .A(n30), .Z(n1685) );
  CIVX2 U1504 ( .A(n87), .Z(n1713) );
  CNIVX1 U1505 ( .A(n116), .Z(n1662) );
  CIVDX2 U1506 ( .A(n55), .Z0(n1567), .Z1(n1568) );
  CIVX2 U1507 ( .A(n1713), .Z(n1712) );
  CNIVX1 U1508 ( .A(n929), .Z(n1570) );
  COR2X1 U1509 ( .A(n723), .B(n738), .Z(n1571) );
  COR2X1 U1510 ( .A(n1574), .B(n630), .Z(n1572) );
  CIVX2 U1511 ( .A(n1709), .Z(n1706) );
  CIVX2 U1512 ( .A(n79), .Z(n1709) );
  COND2X2 U1513 ( .A(n85), .B(n1197), .C(n1196), .D(n82), .Z(n919) );
  CND2X4 U1514 ( .A(n1604), .B(n1605), .Z(n82) );
  CNIVX2 U1515 ( .A(n122), .Z(n1650) );
  CNIVX1 U1516 ( .A(n981), .Z(n1573) );
  COND2XL U1517 ( .A(n112), .B(n1141), .C(n110), .D(n1140), .Z(n868) );
  CIVX3 U1518 ( .A(n1700), .Z(n1699) );
  CND2X2 U1519 ( .A(n95), .B(n1447), .Z(n97) );
  CENX1 U1520 ( .A(n1693), .B(n1651), .Z(n1275) );
  CENX1 U1521 ( .A(n1693), .B(n1653), .Z(n1272) );
  CENXL U1522 ( .A(n1693), .B(n1654), .Z(n1271) );
  CENX1 U1523 ( .A(n1693), .B(n1660), .Z(n1265) );
  CIVX8 U1524 ( .A(n1695), .Z(n1693) );
  CFA1XL U1525 ( .A(n889), .B(n911), .CI(n899), .CO(n508), .S(n509) );
  CENX1 U1526 ( .A(n1714), .B(n1655), .Z(n1162) );
  CIVX2 U1527 ( .A(n1670), .Z(n1668) );
  CIVX4 U1528 ( .A(n1634), .Z(n24) );
  CIVX1 U1529 ( .A(n292), .Z(n291) );
  CIVX2 U1530 ( .A(a[20]), .Z(n1593) );
  CENX1 U1531 ( .A(n1694), .B(n1659), .Z(n1266) );
  CNIVX2 U1532 ( .A(n142), .Z(n1659) );
  COND2XL U1533 ( .A(n77), .B(n1705), .C(n1216), .D(n74), .Z(n857) );
  CENXL U1534 ( .A(n1678), .B(n156), .Z(n1308) );
  CENX1 U1535 ( .A(n1711), .B(n1652), .Z(n1178) );
  CENX2 U1536 ( .A(n1711), .B(a[22]), .Z(n95) );
  CENX1 U1537 ( .A(n1711), .B(n1653), .Z(n1177) );
  COND2X1 U1538 ( .A(n77), .B(n1204), .C(n1203), .D(n74), .Z(n925) );
  COND2XL U1539 ( .A(n61), .B(n1248), .C(n1247), .D(n1639), .Z(n967) );
  CIVX1 U1540 ( .A(n79), .Z(n1710) );
  COND2X1 U1541 ( .A(n107), .B(n1148), .C(n105), .D(n1147), .Z(n874) );
  CEOX2 U1542 ( .A(a[20]), .B(n1712), .Z(n1448) );
  COND2XL U1543 ( .A(n27), .B(n1339), .C(n24), .D(n1338), .Z(n1054) );
  CIVXL U1544 ( .A(n312), .Z(n311) );
  CENX1 U1545 ( .A(n1708), .B(n1651), .Z(n1195) );
  COND2X1 U1546 ( .A(n69), .B(n1232), .C(n1231), .D(n66), .Z(n952) );
  CENX1 U1547 ( .A(n1697), .B(n1650), .Z(n1232) );
  COND2XL U1548 ( .A(n77), .B(n1207), .C(n1206), .D(n74), .Z(n928) );
  CND2IXL U1549 ( .B(n1661), .A(n1706), .Z(n1199) );
  CENXL U1550 ( .A(n1706), .B(n126), .Z(n1194) );
  CND2X2 U1551 ( .A(n1706), .B(a[20]), .Z(n1594) );
  CENXL U1552 ( .A(n1706), .B(n1652), .Z(n1193) );
  CENX2 U1553 ( .A(n1708), .B(n1650), .Z(n1196) );
  CENX1 U1554 ( .A(n1699), .B(n151), .Z(n1217) );
  CFA1XL U1555 ( .A(n989), .B(n1119), .CI(n1035), .CO(n716), .S(n717) );
  CIVX2 U1556 ( .A(n1611), .Z(n262) );
  COND2XL U1557 ( .A(n85), .B(n1709), .C(n1199), .D(n82), .Z(n856) );
  CENX1 U1558 ( .A(n1649), .B(n1716), .Z(n1158) );
  CNIVX2 U1559 ( .A(n130), .Z(n1653) );
  CENX1 U1560 ( .A(n1691), .B(n151), .Z(n1286) );
  CEO3XL U1561 ( .A(n613), .B(n611), .C(n632), .Z(n1574) );
  CNR2IXL U1562 ( .B(n1662), .A(n66), .Z(n955) );
  COND2XL U1563 ( .A(n69), .B(n1220), .C(n1219), .D(n66), .Z(n940) );
  COND2XL U1564 ( .A(n69), .B(n1221), .C(n1220), .D(n66), .Z(n941) );
  CENX1 U1565 ( .A(n1712), .B(n1650), .Z(n1181) );
  COND2X1 U1566 ( .A(n91), .B(n1181), .C(n1180), .D(n89), .Z(n904) );
  CENX1 U1567 ( .A(n1650), .B(n104), .Z(n1148) );
  COND2X1 U1568 ( .A(n61), .B(n1242), .C(n1241), .D(n1639), .Z(n961) );
  CEOX1 U1569 ( .A(a[24]), .B(n1716), .Z(n1446) );
  CIVXL U1570 ( .A(n1710), .Z(n1707) );
  CIVX2 U1571 ( .A(n1710), .Z(n1708) );
  CIVXL U1572 ( .A(n248), .Z(n1575) );
  CENXL U1573 ( .A(n1699), .B(n148), .Z(n1219) );
  CENX1 U1574 ( .A(n1661), .B(n1699), .Z(n1234) );
  COND2X1 U1575 ( .A(n77), .B(n1203), .C(n1202), .D(n74), .Z(n924) );
  CFA1XL U1576 ( .A(n941), .B(n1079), .CI(n1025), .CO(n504), .S(n505) );
  COND2X1 U1577 ( .A(n1159), .B(n102), .C(n100), .D(n1158), .Z(n884) );
  CNR2X1 U1578 ( .A(n234), .B(n239), .Z(n228) );
  CNIVX1 U1579 ( .A(n1030), .Z(n1576) );
  CAN2XL U1580 ( .A(n388), .B(n226), .Z(n1577) );
  COND2X1 U1581 ( .A(n53), .B(n1262), .C(n1261), .D(n50), .Z(n980) );
  COND2X1 U1582 ( .A(n53), .B(n1275), .C(n1274), .D(n50), .Z(n993) );
  CNIVX1 U1583 ( .A(n891), .Z(n1578) );
  CND2X4 U1584 ( .A(n1594), .B(n1595), .Z(n89) );
  CENX1 U1585 ( .A(a[14]), .B(n1699), .Z(n1616) );
  CENXL U1586 ( .A(n1579), .B(n236), .Z(product[26]) );
  CAN2XL U1587 ( .A(n389), .B(n235), .Z(n1579) );
  CENXL U1588 ( .A(n1693), .B(n155), .Z(n1257) );
  CENXL U1589 ( .A(n1686), .B(n155), .Z(n1282) );
  CENXL U1590 ( .A(n1672), .B(n155), .Z(n1338) );
  CIVX3 U1591 ( .A(n1705), .Z(n1701) );
  CNIVX2 U1592 ( .A(n136), .Z(n1656) );
  COND2X1 U1593 ( .A(n27), .B(n1337), .C(n24), .D(n1336), .Z(n1052) );
  COND2X1 U1594 ( .A(n27), .B(n1349), .C(n24), .D(n1348), .Z(n1064) );
  COND2X1 U1595 ( .A(n69), .B(n1226), .C(n1225), .D(n66), .Z(n946) );
  COND2XL U1596 ( .A(n97), .B(n1169), .C(n1168), .D(n95), .Z(n893) );
  COND2XL U1597 ( .A(n97), .B(n1167), .C(n1166), .D(n95), .Z(n891) );
  CENX1 U1598 ( .A(n1664), .B(n153), .Z(n1371) );
  CFA1X1 U1599 ( .A(n924), .B(n1078), .CI(n978), .CO(n478), .S(n479) );
  COND2X1 U1600 ( .A(n53), .B(n1260), .C(n1259), .D(n50), .Z(n978) );
  CEOX1 U1601 ( .A(a[26]), .B(n104), .Z(n1445) );
  CENX1 U1602 ( .A(n1649), .B(n1714), .Z(n1169) );
  CENX1 U1603 ( .A(n1649), .B(n104), .Z(n1149) );
  CANR1X2 U1604 ( .A(n257), .B(n391), .C(n248), .Z(n246) );
  CFA1XL U1605 ( .A(n980), .B(n1080), .CI(n1110), .CO(n528), .S(n529) );
  CFA1XL U1606 ( .A(n940), .B(n1024), .CI(n1050), .CO(n476), .S(n477) );
  CND2X4 U1607 ( .A(n89), .B(n1448), .Z(n91) );
  CENXL U1608 ( .A(n1708), .B(n1660), .Z(n1185) );
  CENXL U1609 ( .A(n1682), .B(n1660), .Z(n1317) );
  CENXL U1610 ( .A(n1671), .B(n1660), .Z(n1346) );
  CENXL U1611 ( .A(n1669), .B(n1660), .Z(n1377) );
  CENXL U1612 ( .A(n1704), .B(n1660), .Z(n1202) );
  CENX1 U1613 ( .A(n1666), .B(n154), .Z(n1370) );
  CENXL U1614 ( .A(n1672), .B(n154), .Z(n1339) );
  CENXL U1615 ( .A(n1679), .B(n154), .Z(n1310) );
  CENXL U1616 ( .A(n1693), .B(n154), .Z(n1258) );
  CND2X1 U1617 ( .A(n391), .B(n1572), .Z(n245) );
  CIVX1 U1618 ( .A(n242), .Z(n241) );
  COND2XL U1619 ( .A(n27), .B(n1333), .C(n24), .D(n1332), .Z(n1048) );
  COND2XL U1620 ( .A(n27), .B(n1334), .C(n24), .D(n1333), .Z(n1049) );
  COND2XL U1621 ( .A(n27), .B(n1356), .C(n24), .D(n1355), .Z(n1071) );
  COND2XL U1622 ( .A(n27), .B(n1358), .C(n24), .D(n1357), .Z(n1073) );
  COND2XL U1623 ( .A(n27), .B(n1354), .C(n24), .D(n1353), .Z(n1069) );
  COND2XL U1624 ( .A(n27), .B(n1350), .C(n24), .D(n1349), .Z(n1065) );
  COND2XL U1625 ( .A(n27), .B(n1357), .C(n24), .D(n1356), .Z(n1072) );
  COND2XL U1626 ( .A(n27), .B(n1353), .C(n24), .D(n1352), .Z(n1068) );
  COND2XL U1627 ( .A(n27), .B(n1335), .C(n24), .D(n1334), .Z(n1050) );
  COND2XL U1628 ( .A(n27), .B(n1341), .C(n24), .D(n1340), .Z(n1056) );
  COND2XL U1629 ( .A(n27), .B(n1347), .C(n24), .D(n1346), .Z(n1062) );
  COND2XL U1630 ( .A(n27), .B(n1355), .C(n24), .D(n1354), .Z(n1070) );
  COND2XL U1631 ( .A(n27), .B(n1338), .C(n24), .D(n1337), .Z(n1053) );
  COND2XL U1632 ( .A(n27), .B(n1351), .C(n24), .D(n1350), .Z(n1066) );
  CNR2IXL U1633 ( .B(n1661), .A(n24), .Z(n1075) );
  COND2XL U1634 ( .A(n27), .B(n1336), .C(n24), .D(n1335), .Z(n1051) );
  COND2XL U1635 ( .A(n27), .B(n1344), .C(n24), .D(n1343), .Z(n1059) );
  COND2XL U1636 ( .A(n27), .B(n1677), .C(n1360), .D(n24), .Z(n863) );
  CENXL U1637 ( .A(n1703), .B(n1659), .Z(n1203) );
  CENXL U1638 ( .A(n1580), .B(n220), .Z(product[28]) );
  CAN2X1 U1639 ( .A(n387), .B(n219), .Z(n1580) );
  CNIVX2 U1640 ( .A(n128), .Z(n1652) );
  CENX1 U1641 ( .A(n1696), .B(n1655), .Z(n1247) );
  COND2X1 U1642 ( .A(n53), .B(n1269), .C(n1268), .D(n50), .Z(n987) );
  CENXL U1643 ( .A(n1712), .B(n1657), .Z(n1173) );
  CENXL U1644 ( .A(n1703), .B(n1657), .Z(n1205) );
  CND2IX4 U1645 ( .B(n1617), .A(n82), .Z(n85) );
  CIVX1 U1646 ( .A(n212), .Z(n210) );
  CNR2IX1 U1647 ( .B(n1661), .A(n105), .Z(n877) );
  COND2XL U1648 ( .A(n36), .B(n1306), .C(n1305), .D(n33), .Z(n1022) );
  COND2XL U1649 ( .A(n36), .B(n1328), .C(n1327), .D(n33), .Z(n1044) );
  COND2XL U1650 ( .A(n36), .B(n1307), .C(n1306), .D(n33), .Z(n1023) );
  COND2XL U1651 ( .A(n36), .B(n1326), .C(n1325), .D(n33), .Z(n1042) );
  COND2XL U1652 ( .A(n36), .B(n1684), .C(n1331), .D(n33), .Z(n862) );
  COND2XL U1653 ( .A(n36), .B(n1318), .C(n1317), .D(n33), .Z(n1034) );
  COND2XL U1654 ( .A(n36), .B(n1323), .C(n1322), .D(n33), .Z(n1039) );
  COND2XL U1655 ( .A(n36), .B(n1309), .C(n1308), .D(n33), .Z(n1025) );
  COND2XL U1656 ( .A(n36), .B(n1330), .C(n1329), .D(n33), .Z(n1046) );
  COND2XL U1657 ( .A(n36), .B(n1319), .C(n1318), .D(n33), .Z(n1035) );
  COND2XL U1658 ( .A(n36), .B(n1308), .C(n1307), .D(n33), .Z(n1024) );
  COND2XL U1659 ( .A(n36), .B(n1329), .C(n1328), .D(n33), .Z(n1045) );
  COND2XL U1660 ( .A(n36), .B(n1314), .C(n1313), .D(n33), .Z(n1030) );
  CNR2IXL U1661 ( .B(n1661), .A(n33), .Z(n1047) );
  CND2IXL U1662 ( .B(n1662), .A(n1568), .Z(n1256) );
  CND2XL U1663 ( .A(n1707), .B(n1649), .Z(n1583) );
  CND2X1 U1664 ( .A(n1581), .B(n1582), .Z(n1584) );
  CND2X1 U1665 ( .A(n1583), .B(n1584), .Z(n1197) );
  CIVXL U1666 ( .A(n1707), .Z(n1581) );
  CIVXL U1667 ( .A(n1649), .Z(n1582) );
  CND2X2 U1668 ( .A(n166), .B(n1586), .Z(n1587) );
  CND2XL U1669 ( .A(n199), .B(n1585), .Z(n1588) );
  CND2X1 U1670 ( .A(n1587), .B(n1588), .Z(product[31]) );
  CIVX2 U1671 ( .A(n166), .Z(n1585) );
  CIVX1 U1672 ( .A(n199), .Z(n1586) );
  COR2XL U1673 ( .A(n107), .B(n1147), .Z(n1589) );
  COR2XL U1674 ( .A(n105), .B(n1146), .Z(n1590) );
  CND2X1 U1675 ( .A(n1589), .B(n1590), .Z(n873) );
  COR2X1 U1676 ( .A(n1569), .B(n1370), .Z(n1592) );
  CND2X2 U1677 ( .A(n1709), .B(n1593), .Z(n1595) );
  COND2XL U1678 ( .A(n91), .B(n1176), .C(n1175), .D(n89), .Z(n899) );
  COND2XL U1679 ( .A(n91), .B(n1180), .C(n1179), .D(n89), .Z(n903) );
  COND2XL U1680 ( .A(n91), .B(n1173), .C(n1172), .D(n89), .Z(n896) );
  COND2X1 U1681 ( .A(n91), .B(n1174), .C(n1173), .D(n89), .Z(n897) );
  COND2X1 U1682 ( .A(n91), .B(n1175), .C(n1174), .D(n89), .Z(n898) );
  CNR2XL U1683 ( .A(n1246), .B(n1639), .Z(n1597) );
  COR2X1 U1684 ( .A(n1596), .B(n1597), .Z(n966) );
  CND2X4 U1685 ( .A(n1452), .B(n1638), .Z(n61) );
  CND2XL U1686 ( .A(n1703), .B(n1654), .Z(n1600) );
  CND2X1 U1687 ( .A(n1598), .B(n1599), .Z(n1601) );
  CND2X1 U1688 ( .A(n1600), .B(n1601), .Z(n1208) );
  CIVX1 U1689 ( .A(n1703), .Z(n1598) );
  CIVXL U1690 ( .A(n1654), .Z(n1599) );
  CIVXL U1691 ( .A(n1705), .Z(n1703) );
  CNIVX4 U1692 ( .A(n132), .Z(n1654) );
  CND2X1 U1693 ( .A(n1701), .B(a[18]), .Z(n1604) );
  CND2X1 U1694 ( .A(n1602), .B(n1603), .Z(n1605) );
  CIVX2 U1695 ( .A(n1701), .Z(n1602) );
  CIVX2 U1696 ( .A(a[18]), .Z(n1603) );
  COND2XL U1697 ( .A(n85), .B(n1189), .C(n1188), .D(n82), .Z(n911) );
  COND2XL U1698 ( .A(n85), .B(n1187), .C(n1186), .D(n82), .Z(n909) );
  COND2XL U1699 ( .A(n85), .B(n1186), .C(n1185), .D(n82), .Z(n908) );
  CND2X1 U1700 ( .A(a[22]), .B(n1607), .Z(n1608) );
  CND2X1 U1701 ( .A(n1606), .B(n1714), .Z(n1609) );
  CIVXL U1702 ( .A(a[22]), .Z(n1606) );
  CIVX2 U1703 ( .A(n1714), .Z(n1607) );
  CENXL U1704 ( .A(n1666), .B(n1653), .Z(n1384) );
  CENXL U1705 ( .A(n1706), .B(n1653), .Z(n1192) );
  CENXL U1706 ( .A(n1714), .B(n1653), .Z(n1164) );
  COND2XL U1707 ( .A(n107), .B(n1146), .C(n105), .D(n1145), .Z(n872) );
  COND2XL U1708 ( .A(n107), .B(n1470), .C(n105), .D(n1151), .Z(n852) );
  CENXL U1709 ( .A(n1712), .B(n1655), .Z(n1175) );
  COND2XL U1710 ( .A(n102), .B(n1717), .C(n100), .D(n1160), .Z(n853) );
  CENX2 U1711 ( .A(n1714), .B(a[24]), .Z(n100) );
  CENXL U1712 ( .A(n1661), .B(n113), .Z(n1138) );
  CENXL U1713 ( .A(n1681), .B(n1661), .Z(n1330) );
  CENXL U1714 ( .A(n1661), .B(n109), .Z(n1143) );
  CENXL U1715 ( .A(n1661), .B(n1568), .Z(n1255) );
  CENXL U1716 ( .A(n1661), .B(n1707), .Z(n1198) );
  CENXL U1717 ( .A(n1661), .B(n1694), .Z(n1278) );
  CENXL U1718 ( .A(n1661), .B(n104), .Z(n1150) );
  CENXL U1719 ( .A(n1661), .B(n1703), .Z(n1215) );
  CENXL U1720 ( .A(n1661), .B(n1712), .Z(n1183) );
  CENXL U1721 ( .A(n1661), .B(n1716), .Z(n1159) );
  CENXL U1722 ( .A(n1661), .B(n1714), .Z(n1170) );
  CENXL U1723 ( .A(n1714), .B(n1656), .Z(n1161) );
  CENXL U1724 ( .A(n1675), .B(n1656), .Z(n1350) );
  CENXL U1725 ( .A(n1689), .B(n1656), .Z(n1294) );
  CENXL U1726 ( .A(n1669), .B(n1656), .Z(n1381) );
  CENXL U1727 ( .A(n1681), .B(n1656), .Z(n1321) );
  CENXL U1728 ( .A(n1694), .B(n1656), .Z(n1269) );
  CENXL U1729 ( .A(n1707), .B(n1656), .Z(n1189) );
  CENXL U1730 ( .A(n1696), .B(n1656), .Z(n1246) );
  CENXL U1731 ( .A(n1712), .B(n1656), .Z(n1174) );
  CENXL U1732 ( .A(n1698), .B(n150), .Z(n1218) );
  CENXL U1733 ( .A(n1568), .B(n150), .Z(n1239) );
  CENXL U1734 ( .A(n1664), .B(n150), .Z(n1374) );
  CENXL U1735 ( .A(n1671), .B(n150), .Z(n1343) );
  CENXL U1736 ( .A(n1683), .B(n150), .Z(n1314) );
  CENXL U1737 ( .A(n1694), .B(n150), .Z(n1262) );
  CHA1XL U1738 ( .A(n854), .B(n904), .CO(n628), .S(n629) );
  CENXL U1739 ( .A(n1714), .B(n126), .Z(n1166) );
  CENXL U1740 ( .A(n1714), .B(n1651), .Z(n1167) );
  CENXL U1741 ( .A(n1668), .B(b[29]), .Z(n1361) );
  CENXL U1742 ( .A(n1668), .B(n1661), .Z(n1390) );
  CEOX2 U1743 ( .A(n1668), .B(a[4]), .Z(n1634) );
  CENXL U1744 ( .A(n1714), .B(n1650), .Z(n1168) );
  CANR1X1 U1745 ( .A(n1619), .B(n213), .C(n1618), .Z(n199) );
  CENXL U1746 ( .A(n1712), .B(n1649), .Z(n1182) );
  CENXL U1747 ( .A(n1668), .B(n1649), .Z(n1389) );
  CND2X1 U1748 ( .A(n631), .B(n650), .Z(n270) );
  CENXL U1749 ( .A(n1648), .B(n208), .Z(product[30]) );
  CND2X1 U1750 ( .A(n1699), .B(a[16]), .Z(n1613) );
  CND2X2 U1751 ( .A(n1700), .B(n1612), .Z(n1614) );
  CND2X4 U1752 ( .A(n1613), .B(n1614), .Z(n74) );
  CNR2X1 U1753 ( .A(n245), .B(n261), .Z(n243) );
  CENX1 U1754 ( .A(n1689), .B(n146), .Z(n1289) );
  CENX1 U1755 ( .A(n1682), .B(n146), .Z(n1316) );
  CENX1 U1756 ( .A(n1671), .B(n146), .Z(n1345) );
  CENX1 U1757 ( .A(n1694), .B(n146), .Z(n1264) );
  COND1X1 U1758 ( .A(n352), .B(n340), .C(n341), .Z(n339) );
  CIVX1 U1759 ( .A(n21), .Z(n1677) );
  CANR1X2 U1760 ( .A(n308), .B(n1571), .C(n301), .Z(n299) );
  CND2X1 U1761 ( .A(n819), .B(n826), .Z(n350) );
  COND1XL U1762 ( .A(n368), .B(n366), .C(n367), .Z(n365) );
  COR2X1 U1763 ( .A(n847), .B(n848), .Z(n1630) );
  CEO3X1 U1764 ( .A(n434), .B(n416), .C(n432), .Z(n415) );
  CEO3X1 U1765 ( .A(n436), .B(n418), .C(n417), .Z(n416) );
  CENX1 U1766 ( .A(n1666), .B(n1654), .Z(n1383) );
  CNR2IXL U1767 ( .B(n1661), .A(n89), .Z(n907) );
  CNIVX1 U1768 ( .A(n144), .Z(n1660) );
  CEOX2 U1769 ( .A(n1675), .B(a[6]), .Z(n1633) );
  COND1X1 U1770 ( .A(n214), .B(n1559), .C(n215), .Z(n213) );
  CANR1X1 U1771 ( .A(n229), .B(n216), .C(n217), .Z(n215) );
  CEOXL U1772 ( .A(n176), .B(n278), .Z(product[21]) );
  CND2XL U1773 ( .A(n394), .B(n1640), .Z(n176) );
  CEOXL U1774 ( .A(n1615), .B(n213), .Z(product[29]) );
  CAN2XL U1775 ( .A(n1620), .B(n212), .Z(n1615) );
  CND2XL U1776 ( .A(n390), .B(n240), .Z(n172) );
  CND2XL U1777 ( .A(n320), .B(n1624), .Z(n313) );
  CIVX1 U1778 ( .A(n318), .Z(n316) );
  CEOXL U1779 ( .A(n177), .B(n286), .Z(product[20]) );
  CND2XL U1780 ( .A(n395), .B(n285), .Z(n177) );
  CEOXL U1781 ( .A(n183), .B(n324), .Z(product[14]) );
  CND2XL U1782 ( .A(n401), .B(n323), .Z(n183) );
  CEOXL U1783 ( .A(n182), .B(n319), .Z(product[15]) );
  CND2XL U1784 ( .A(n1624), .B(n318), .Z(n182) );
  CEOXL U1785 ( .A(n181), .B(n311), .Z(product[16]) );
  CND2X1 U1786 ( .A(n1571), .B(n399), .Z(n298) );
  CND2XL U1787 ( .A(n1625), .B(n290), .Z(n178) );
  COR2XL U1788 ( .A(n459), .B(n486), .Z(n1620) );
  CNIVXL U1789 ( .A(n273), .Z(n1640) );
  CND2XL U1790 ( .A(n1627), .B(n1626), .Z(n340) );
  CNR2X1 U1791 ( .A(n739), .B(n752), .Z(n305) );
  CND2XL U1792 ( .A(n1627), .B(n345), .Z(n187) );
  CND2XL U1793 ( .A(n404), .B(n337), .Z(n186) );
  CEOXL U1794 ( .A(n186), .B(n338), .Z(product[11]) );
  CND2XL U1795 ( .A(n671), .B(n688), .Z(n285) );
  CND2XL U1796 ( .A(n1628), .B(n356), .Z(n189) );
  CND2XL U1797 ( .A(n1626), .B(n350), .Z(n188) );
  CND2XL U1798 ( .A(n402), .B(n328), .Z(n184) );
  CND2XL U1799 ( .A(n430), .B(n415), .Z(n198) );
  CND2XL U1800 ( .A(n408), .B(n359), .Z(n190) );
  CEOXL U1801 ( .A(n360), .B(n190), .Z(product[7]) );
  CND2XL U1802 ( .A(n1631), .B(n364), .Z(n191) );
  CND2XL U1803 ( .A(n843), .B(n846), .Z(n367) );
  CND2XL U1804 ( .A(n849), .B(n864), .Z(n375) );
  CANR1X1 U1805 ( .A(n373), .B(n1630), .C(n370), .Z(n368) );
  CND2XL U1806 ( .A(n1630), .B(n372), .Z(n193) );
  COR2XL U1807 ( .A(n1135), .B(n1105), .Z(n1632) );
  CIVX3 U1808 ( .A(n1636), .Z(n1639) );
  CIVX3 U1809 ( .A(n1717), .Z(n1716) );
  CIVX3 U1810 ( .A(n1692), .Z(n1688) );
  CNR2IXL U1811 ( .B(n1662), .A(n1569), .Z(n1105) );
  COND2XL U1812 ( .A(n27), .B(n1359), .C(n24), .D(n1358), .Z(n1074) );
  CND2XL U1813 ( .A(n412), .B(n375), .Z(n194) );
  CEOXL U1814 ( .A(n376), .B(n194), .Z(product[3]) );
  CENX4 U1815 ( .A(n1696), .B(a[14]), .Z(n66) );
  CND2X2 U1816 ( .A(n100), .B(n1446), .Z(n102) );
  CND2IX4 U1817 ( .B(n1616), .A(n66), .Z(n69) );
  CENXL U1818 ( .A(n1690), .B(n150), .Z(n1287) );
  CND2XL U1819 ( .A(n1443), .B(n114), .Z(n115) );
  CEOXL U1820 ( .A(a[30]), .B(n113), .Z(n1443) );
  CND2XL U1821 ( .A(n1632), .B(n380), .Z(n195) );
  CANR1XL U1822 ( .A(n390), .B(n241), .C(n238), .Z(n236) );
  CENX1 U1823 ( .A(n260), .B(n174), .Z(product[23]) );
  CND2XL U1824 ( .A(n1572), .B(n259), .Z(n174) );
  CANR1XL U1825 ( .A(n1620), .B(n213), .C(n210), .Z(n208) );
  COND1XL U1826 ( .A(n223), .B(n231), .C(n226), .Z(n222) );
  CNR2IXL U1827 ( .B(n228), .A(n223), .Z(n221) );
  CANR1XL U1828 ( .A(n1572), .B(n1611), .C(n257), .Z(n253) );
  CENX1 U1829 ( .A(n251), .B(n173), .Z(product[24]) );
  CND2XL U1830 ( .A(n391), .B(n1575), .Z(n173) );
  COND1XL U1831 ( .A(n252), .B(n278), .C(n253), .Z(n251) );
  CND2XL U1832 ( .A(n263), .B(n1572), .Z(n252) );
  CANR1XL U1833 ( .A(n221), .B(n241), .C(n222), .Z(n220) );
  CAOR1X1 U1834 ( .A(n210), .B(n1621), .C(n205), .Z(n1618) );
  CNR2XL U1835 ( .A(n295), .B(n298), .Z(n293) );
  CND2X1 U1836 ( .A(n395), .B(n1625), .Z(n280) );
  CNR2X1 U1837 ( .A(n487), .B(n512), .Z(n218) );
  CNR2X1 U1838 ( .A(n513), .B(n538), .Z(n223) );
  CENX1 U1839 ( .A(n297), .B(n179), .Z(product[18]) );
  CND2X1 U1840 ( .A(n397), .B(n296), .Z(n179) );
  CENX1 U1841 ( .A(n271), .B(n175), .Z(product[22]) );
  CND2XL U1842 ( .A(n393), .B(n270), .Z(n175) );
  COND1XL U1843 ( .A(n272), .B(n278), .C(n1640), .Z(n271) );
  CENX1 U1844 ( .A(n304), .B(n180), .Z(product[17]) );
  CND2XL U1845 ( .A(n1571), .B(n303), .Z(n180) );
  COND1XL U1846 ( .A(n305), .B(n311), .C(n306), .Z(n304) );
  CENX1 U1847 ( .A(n291), .B(n178), .Z(product[19]) );
  CANR1XL U1848 ( .A(n1625), .B(n291), .C(n288), .Z(n286) );
  CANR1XL U1849 ( .A(n402), .B(n329), .C(n326), .Z(n324) );
  CANR1XL U1850 ( .A(n320), .B(n329), .C(n321), .Z(n319) );
  CND2XL U1851 ( .A(n399), .B(n306), .Z(n181) );
  CND2X1 U1852 ( .A(n563), .B(n586), .Z(n240) );
  CND2X1 U1853 ( .A(n393), .B(n394), .Z(n261) );
  COR2X1 U1854 ( .A(n431), .B(n458), .Z(n1621) );
  CND2X1 U1855 ( .A(n459), .B(n486), .Z(n212) );
  CND2X1 U1856 ( .A(n487), .B(n512), .Z(n219) );
  CND2X1 U1857 ( .A(n431), .B(n458), .Z(n207) );
  CANR1XL U1858 ( .A(n348), .B(n1627), .C(n343), .Z(n341) );
  CENX1 U1859 ( .A(n1622), .B(n633), .Z(n631) );
  CENX1 U1860 ( .A(n635), .B(n652), .Z(n1622) );
  CENX1 U1861 ( .A(n1623), .B(n489), .Z(n487) );
  CENX1 U1862 ( .A(n514), .B(n491), .Z(n1623) );
  CNR2XL U1863 ( .A(n333), .B(n336), .Z(n331) );
  CENX1 U1864 ( .A(n188), .B(n351), .Z(product[9]) );
  CENX1 U1865 ( .A(n335), .B(n185), .Z(product[12]) );
  CND2X1 U1866 ( .A(n403), .B(n334), .Z(n185) );
  COND1XL U1867 ( .A(n336), .B(n338), .C(n337), .Z(n335) );
  CENX1 U1868 ( .A(n329), .B(n184), .Z(product[13]) );
  CNR2X1 U1869 ( .A(n322), .B(n327), .Z(n320) );
  CNR2X1 U1870 ( .A(n671), .B(n688), .Z(n284) );
  CEOX1 U1871 ( .A(n346), .B(n187), .Z(product[10]) );
  CANR1XL U1872 ( .A(n1626), .B(n351), .C(n348), .Z(n346) );
  COR2X1 U1873 ( .A(n753), .B(n766), .Z(n1624) );
  COR2X1 U1874 ( .A(n689), .B(n706), .Z(n1625) );
  CND2X1 U1875 ( .A(n689), .B(n706), .Z(n290) );
  CND2X1 U1876 ( .A(n707), .B(n722), .Z(n296) );
  CND2X1 U1877 ( .A(n753), .B(n766), .Z(n318) );
  CND2X1 U1878 ( .A(n767), .B(n778), .Z(n323) );
  CENX1 U1879 ( .A(n189), .B(n357), .Z(product[8]) );
  CANR1XL U1880 ( .A(n365), .B(n1631), .C(n362), .Z(n360) );
  CNR2X1 U1881 ( .A(n801), .B(n810), .Z(n336) );
  CNR2X1 U1882 ( .A(n779), .B(n790), .Z(n327) );
  CND2X1 U1883 ( .A(n1629), .B(n198), .Z(n166) );
  COR2X1 U1884 ( .A(n819), .B(n826), .Z(n1626) );
  COR2X1 U1885 ( .A(n811), .B(n818), .Z(n1627) );
  CND2X1 U1886 ( .A(n801), .B(n810), .Z(n337) );
  CND2X1 U1887 ( .A(n827), .B(n832), .Z(n356) );
  CND2X1 U1888 ( .A(n811), .B(n818), .Z(n345) );
  CND2X1 U1889 ( .A(n791), .B(n800), .Z(n334) );
  COR2X1 U1890 ( .A(n827), .B(n832), .Z(n1628) );
  COR2X1 U1891 ( .A(n430), .B(n415), .Z(n1629) );
  CENX1 U1892 ( .A(n191), .B(n365), .Z(product[6]) );
  CEOX1 U1893 ( .A(n368), .B(n192), .Z(product[5]) );
  CND2X1 U1894 ( .A(n410), .B(n367), .Z(n192) );
  CNR2X1 U1895 ( .A(n833), .B(n838), .Z(n358) );
  CNR2X1 U1896 ( .A(n843), .B(n846), .Z(n366) );
  CNR2X1 U1897 ( .A(n849), .B(n864), .Z(n374) );
  CND2X1 U1898 ( .A(n833), .B(n838), .Z(n359) );
  CND2X1 U1899 ( .A(n847), .B(n848), .Z(n372) );
  CND2X1 U1900 ( .A(n839), .B(n842), .Z(n364) );
  CND2X1 U1901 ( .A(n1135), .B(n1105), .Z(n380) );
  COR2X1 U1902 ( .A(n839), .B(n842), .Z(n1631) );
  CENX1 U1903 ( .A(n193), .B(n373), .Z(product[4]) );
  COND1XL U1904 ( .A(n376), .B(n374), .C(n375), .Z(n373) );
  CENX1 U1905 ( .A(n1694), .B(n1658), .Z(n1267) );
  CENX1 U1906 ( .A(n1697), .B(n1651), .Z(n1231) );
  CENX1 U1907 ( .A(n1679), .B(n1654), .Z(n1323) );
  CENX1 U1908 ( .A(n1698), .B(n1658), .Z(n1223) );
  CENX1 U1909 ( .A(n1671), .B(n1658), .Z(n1348) );
  CENX1 U1910 ( .A(n1675), .B(n1661), .Z(n1359) );
  CENX1 U1911 ( .A(n1654), .B(n1716), .Z(n1152) );
  CENX1 U1912 ( .A(n1712), .B(n1658), .Z(n1172) );
  CENX1 U1913 ( .A(n1698), .B(n1652), .Z(n1229) );
  CNR2IX1 U1914 ( .B(n1661), .A(n100), .Z(n885) );
  CENX1 U1915 ( .A(n1669), .B(n1658), .Z(n1379) );
  CENX1 U1916 ( .A(n1690), .B(n1660), .Z(n1290) );
  CENX1 U1917 ( .A(n1712), .B(n1651), .Z(n1180) );
  CENX1 U1918 ( .A(n1689), .B(n1658), .Z(n1292) );
  CENX1 U1919 ( .A(n1708), .B(n1654), .Z(n1191) );
  CENX1 U1920 ( .A(n1687), .B(n1651), .Z(n1300) );
  CENX1 U1921 ( .A(n1681), .B(n1655), .Z(n1322) );
  CENX1 U1922 ( .A(n1681), .B(n1658), .Z(n1319) );
  CENX1 U1923 ( .A(n1688), .B(n1655), .Z(n1295) );
  CENX1 U1924 ( .A(n1708), .B(n1655), .Z(n1190) );
  CENX1 U1925 ( .A(n1712), .B(n1654), .Z(n1176) );
  CENX1 U1926 ( .A(n1708), .B(n1658), .Z(n1187) );
  CENX1 U1927 ( .A(n1652), .B(n1716), .Z(n1154) );
  CENXL U1928 ( .A(n1674), .B(n1657), .Z(n1349) );
  CENX1 U1929 ( .A(n1714), .B(n1652), .Z(n1165) );
  CENX1 U1930 ( .A(n1693), .B(n1652), .Z(n1273) );
  CENX1 U1931 ( .A(n1669), .B(n1655), .Z(n1382) );
  CENX1 U1932 ( .A(n1687), .B(n1661), .Z(n1303) );
  CENX1 U1933 ( .A(n1714), .B(n1654), .Z(n1163) );
  CENX1 U1934 ( .A(n1667), .B(n1651), .Z(n1387) );
  CENX1 U1935 ( .A(n1667), .B(n1652), .Z(n1385) );
  CNR2IX1 U1936 ( .B(n1661), .A(n110), .Z(n871) );
  CNR2IXL U1937 ( .B(n1662), .A(n1639), .Z(n975) );
  CNR2IX1 U1938 ( .B(n1661), .A(n82), .Z(n921) );
  CNR2IX1 U1939 ( .B(n1661), .A(n114), .Z(n867) );
  CNR2IX1 U1940 ( .B(n1661), .A(n42), .Z(n1021) );
  CNIVX1 U1941 ( .A(n930), .Z(n1641) );
  CEOX1 U1942 ( .A(n872), .B(n850), .Z(n429) );
  CNR2IX1 U1943 ( .B(n1662), .A(n1564), .Z(product[0]) );
  CENX1 U1944 ( .A(n1690), .B(n148), .Z(n1288) );
  CENX1 U1945 ( .A(n1683), .B(n152), .Z(n1312) );
  CENX1 U1946 ( .A(n1697), .B(n146), .Z(n1220) );
  CENX1 U1947 ( .A(n1686), .B(n156), .Z(n1281) );
  CENX1 U1948 ( .A(n1652), .B(n104), .Z(n1145) );
  CENX1 U1949 ( .A(n104), .B(a[28]), .Z(n110) );
  CENX1 U1950 ( .A(n1688), .B(n157), .Z(n1280) );
  CENX1 U1951 ( .A(n1665), .B(n148), .Z(n1375) );
  CENX1 U1952 ( .A(n109), .B(a[30]), .Z(n114) );
  CENX1 U1953 ( .A(n1669), .B(n146), .Z(n1376) );
  CENX1 U1954 ( .A(n1694), .B(n151), .Z(n1261) );
  CENX1 U1955 ( .A(n1694), .B(n152), .Z(n1260) );
  CENX1 U1956 ( .A(n1704), .B(n146), .Z(n1201) );
  CIVX4 U1957 ( .A(n1633), .Z(n33) );
  CENX1 U1958 ( .A(n1651), .B(n109), .Z(n1140) );
  CENX1 U1959 ( .A(n1690), .B(n152), .Z(n1285) );
  CENX1 U1960 ( .A(n1678), .B(n153), .Z(n1311) );
  CENX1 U1961 ( .A(n1678), .B(n157), .Z(n1307) );
  CENX1 U1962 ( .A(n1678), .B(b[24]), .Z(n1306) );
  CENX1 U1963 ( .A(n1665), .B(n157), .Z(n1367) );
  CENX1 U1964 ( .A(n1665), .B(n156), .Z(n1368) );
  CENX1 U1965 ( .A(n1671), .B(b[24]), .Z(n1335) );
  CENX1 U1966 ( .A(n1671), .B(b[25]), .Z(n1334) );
  CENX1 U1967 ( .A(n1671), .B(b[26]), .Z(n1333) );
  CIVX2 U1968 ( .A(n1636), .Z(n1638) );
  CENX1 U1969 ( .A(n1665), .B(b[24]), .Z(n1366) );
  CENX1 U1970 ( .A(n1704), .B(n148), .Z(n1200) );
  CENX1 U1971 ( .A(n1665), .B(b[25]), .Z(n1365) );
  CENX1 U1972 ( .A(n1664), .B(b[26]), .Z(n1364) );
  CENX1 U1973 ( .A(n1664), .B(b[27]), .Z(n1363) );
  CENX1 U1974 ( .A(n1664), .B(b[28]), .Z(n1362) );
  CND2X1 U1975 ( .A(n1444), .B(n110), .Z(n112) );
  CEOX1 U1976 ( .A(a[28]), .B(n109), .Z(n1444) );
  CEOX2 U1977 ( .A(n1693), .B(a[12]), .Z(n1636) );
  CIVX2 U1979 ( .A(n71), .Z(n1705) );
  CIVX2 U1980 ( .A(n1670), .Z(n1667) );
  CIVX3 U1981 ( .A(n12), .Z(n1670) );
  COND2XL U1982 ( .A(n53), .B(n1258), .C(n1257), .D(n50), .Z(n976) );
  COND2XL U1983 ( .A(n53), .B(n1259), .C(n1258), .D(n50), .Z(n977) );
  COND2XL U1984 ( .A(n53), .B(n1274), .C(n1273), .D(n50), .Z(n992) );
  CNR2IXL U1985 ( .B(n1662), .A(n50), .Z(n997) );
  COND2XL U1986 ( .A(n53), .B(n1272), .C(n1271), .D(n50), .Z(n990) );
  COND2XL U1987 ( .A(n53), .B(n1270), .C(n1269), .D(n50), .Z(n988) );
  COND2XL U1988 ( .A(n53), .B(n1278), .C(n1277), .D(n50), .Z(n996) );
  COND2XL U1989 ( .A(n53), .B(n1266), .C(n1265), .D(n50), .Z(n984) );
  COND2XL U1990 ( .A(n53), .B(n1265), .C(n1264), .D(n50), .Z(n983) );
  COND2XL U1991 ( .A(n53), .B(n1271), .C(n1270), .D(n50), .Z(n989) );
  COND2XL U1992 ( .A(n53), .B(n1263), .C(n1262), .D(n50), .Z(n981) );
  COND2XL U1993 ( .A(n53), .B(n1276), .C(n1275), .D(n50), .Z(n994) );
  COND2XL U1994 ( .A(n53), .B(n1277), .C(n1276), .D(n50), .Z(n995) );
  COND2XL U1995 ( .A(n53), .B(n1264), .C(n1263), .D(n50), .Z(n982) );
  CIVX1 U1996 ( .A(n1677), .Z(n1676) );
  CENX1 U1997 ( .A(a[6]), .B(n1684), .Z(n1455) );
  CIVX3 U1998 ( .A(n48), .Z(n1695) );
  CIVX2 U1999 ( .A(n1692), .Z(n1691) );
  CIVX1 U2000 ( .A(n1700), .Z(n1697) );
  CNR2X1 U2001 ( .A(n563), .B(n586), .Z(n239) );
  COAN1X1 U2002 ( .A(n290), .B(n284), .C(n285), .Z(n281) );
  CNR2X1 U2003 ( .A(n651), .B(n670), .Z(n272) );
  COND2XL U2004 ( .A(n53), .B(n1695), .C(n1279), .D(n50), .Z(n860) );
  CND2IXL U2005 ( .B(n1661), .A(n1694), .Z(n1279) );
  CFA1XL U2006 ( .A(n1041), .B(n1095), .CI(n1067), .CO(n796), .S(n797) );
  COND2XL U2007 ( .A(n61), .B(n1567), .C(n1256), .D(n1639), .Z(n859) );
  CIVX1 U2008 ( .A(n1670), .Z(n1669) );
  CND2XL U2009 ( .A(n489), .B(n491), .Z(n1642) );
  CND2XL U2010 ( .A(n489), .B(n514), .Z(n1643) );
  CND2XL U2011 ( .A(n491), .B(n514), .Z(n1644) );
  CND3XL U2012 ( .A(n1642), .B(n1643), .C(n1644), .Z(n486) );
  CFA1XL U2013 ( .A(n928), .B(n1082), .CI(n982), .CO(n580), .S(n581) );
  COND2XL U2014 ( .A(n27), .B(n1340), .C(n24), .D(n1339), .Z(n1055) );
  CIVX1 U2015 ( .A(n1677), .Z(n1671) );
  CIVX1 U2016 ( .A(n1692), .Z(n1690) );
  COND2XL U2017 ( .A(n18), .B(n1366), .C(n1569), .D(n1365), .Z(n1080) );
  CIVX1 U2018 ( .A(n1670), .Z(n1665) );
  CENX1 U2019 ( .A(n1666), .B(n155), .Z(n1369) );
  COND2XL U2020 ( .A(n69), .B(n1700), .C(n1235), .D(n66), .Z(n858) );
  COND2XL U2021 ( .A(n69), .B(n1219), .C(n1218), .D(n66), .Z(n939) );
  COND2XL U2022 ( .A(n69), .B(n1218), .C(n1217), .D(n66), .Z(n938) );
  COND2XL U2023 ( .A(n69), .B(n1230), .C(n1229), .D(n66), .Z(n950) );
  CIVX2 U2024 ( .A(n1713), .Z(n1711) );
  COND2XL U2025 ( .A(n27), .B(n1352), .C(n24), .D(n1351), .Z(n1067) );
  CENX1 U2026 ( .A(n1673), .B(n1654), .Z(n1352) );
  CENX1 U2027 ( .A(n1673), .B(n1652), .Z(n1354) );
  CENX1 U2028 ( .A(n1676), .B(n152), .Z(n1341) );
  CIVX1 U2029 ( .A(n239), .Z(n390) );
  CND2X1 U2030 ( .A(n513), .B(n538), .Z(n226) );
  CND2X1 U2031 ( .A(n539), .B(n562), .Z(n235) );
  CIVXL U2032 ( .A(n223), .Z(n388) );
  COND2XL U2033 ( .A(n18), .B(n1362), .C(n1569), .D(n1361), .Z(n1076) );
  COND2XL U2034 ( .A(n18), .B(n1363), .C(n1569), .D(n1362), .Z(n1077) );
  COND2XL U2035 ( .A(n18), .B(n1670), .C(n1391), .D(n1569), .Z(n864) );
  COND2XL U2036 ( .A(n18), .B(n1388), .C(n1569), .D(n1387), .Z(n1102) );
  COND2XL U2037 ( .A(n18), .B(n1385), .C(n1569), .D(n1384), .Z(n1099) );
  COND2XL U2038 ( .A(n18), .B(n1383), .C(n1569), .D(n1382), .Z(n1097) );
  COND2XL U2039 ( .A(n18), .B(n1386), .C(n1569), .D(n1385), .Z(n1100) );
  COND2XL U2040 ( .A(n18), .B(n1384), .C(n1569), .D(n1383), .Z(n1098) );
  COND2XL U2041 ( .A(n18), .B(n1390), .C(n1569), .D(n1389), .Z(n1104) );
  COND2XL U2042 ( .A(n18), .B(n1365), .C(n1569), .D(n1364), .Z(n1079) );
  COND2XL U2043 ( .A(n18), .B(n1364), .C(n1569), .D(n1363), .Z(n1078) );
  COND2XL U2044 ( .A(n18), .B(n1389), .C(n1569), .D(n1388), .Z(n1103) );
  COND2XL U2045 ( .A(n18), .B(n1370), .C(n1569), .D(n1369), .Z(n1084) );
  COND2XL U2046 ( .A(n18), .B(n1376), .C(n1569), .D(n1375), .Z(n1090) );
  COND2XL U2047 ( .A(n18), .B(n1387), .C(n1569), .D(n1386), .Z(n1101) );
  COND2XL U2048 ( .A(n18), .B(n1378), .C(n1569), .D(n1377), .Z(n1092) );
  CENX1 U2049 ( .A(n1672), .B(n156), .Z(n1337) );
  CENX1 U2050 ( .A(n1672), .B(n157), .Z(n1336) );
  CIVX3 U2051 ( .A(n1695), .Z(n1694) );
  CIVX1 U2052 ( .A(n1685), .Z(n1681) );
  COND2XL U2053 ( .A(n36), .B(n1325), .C(n1324), .D(n33), .Z(n1041) );
  CENX1 U2054 ( .A(n1680), .B(n1652), .Z(n1325) );
  CENX1 U2055 ( .A(n1680), .B(n1651), .Z(n1327) );
  CIVXL U2056 ( .A(n229), .Z(n231) );
  CIVX1 U2057 ( .A(n1692), .Z(n1687) );
  CANR1X2 U2058 ( .A(n331), .B(n339), .C(n332), .Z(n330) );
  CIVXL U2059 ( .A(n1705), .Z(n1704) );
  CENX1 U2060 ( .A(n1563), .B(n1651), .Z(n1212) );
  CEOX1 U2061 ( .A(a[16]), .B(n1701), .Z(n1450) );
  CND2IXL U2062 ( .B(n1661), .A(n1701), .Z(n1216) );
  CENX1 U2063 ( .A(n1704), .B(n1658), .Z(n1204) );
  CFA1X1 U2064 ( .A(n900), .B(n960), .CI(n926), .CO(n532), .S(n533) );
  COND2X1 U2065 ( .A(n77), .B(n1205), .C(n1204), .D(n74), .Z(n926) );
  CIVXL U2066 ( .A(n234), .Z(n389) );
  COND2XL U2067 ( .A(n44), .B(n1692), .C(n1304), .D(n42), .Z(n861) );
  CND2IXL U2068 ( .B(n1662), .A(n1686), .Z(n1304) );
  CENX1 U2069 ( .A(n1686), .B(n154), .Z(n1283) );
  CENX1 U2070 ( .A(n1686), .B(n153), .Z(n1284) );
  CIVX1 U2071 ( .A(n1670), .Z(n1664) );
  CIVX2 U2072 ( .A(n1684), .Z(n1678) );
  CFA1X1 U2073 ( .A(n921), .B(n951), .CI(n935), .CO(n720), .S(n721) );
  COND2X1 U2074 ( .A(n77), .B(n1214), .C(n1213), .D(n74), .Z(n935) );
  CENXL U2075 ( .A(n1679), .B(n1653), .Z(n1324) );
  CENX1 U2076 ( .A(n1679), .B(n155), .Z(n1309) );
  CFA1X1 U2077 ( .A(n931), .B(n1057), .CI(n985), .CO(n646), .S(n647) );
  COND2X1 U2078 ( .A(n77), .B(n1210), .C(n1209), .D(n74), .Z(n931) );
  CENX1 U2079 ( .A(n1687), .B(n1654), .Z(n1296) );
  CIVX1 U2080 ( .A(n1692), .Z(n1689) );
  CND2X1 U2081 ( .A(n216), .B(n228), .Z(n214) );
  COND2X1 U2082 ( .A(n77), .B(n1211), .C(n1210), .D(n74), .Z(n932) );
  CENX1 U2083 ( .A(n1698), .B(n1656), .Z(n1225) );
  CENX1 U2084 ( .A(n1698), .B(n1654), .Z(n1227) );
  COND2X1 U2085 ( .A(n77), .B(n1213), .C(n1212), .D(n74), .Z(n934) );
  COND1XL U2086 ( .A(n298), .B(n311), .C(n299), .Z(n297) );
  CND2XL U2087 ( .A(n633), .B(n652), .Z(n1645) );
  CND2X1 U2088 ( .A(n633), .B(n635), .Z(n1646) );
  CND2XL U2089 ( .A(n652), .B(n635), .Z(n1647) );
  CNR2X1 U2090 ( .A(n218), .B(n223), .Z(n216) );
  COND2XL U2091 ( .A(n97), .B(n1162), .C(n1161), .D(n95), .Z(n886) );
  COND2XL U2092 ( .A(n97), .B(n1164), .C(n1163), .D(n95), .Z(n888) );
  COND2XL U2093 ( .A(n97), .B(n1168), .C(n1167), .D(n95), .Z(n892) );
  COND2XL U2094 ( .A(n97), .B(n1715), .C(n95), .D(n1171), .Z(n854) );
  CND2IXL U2095 ( .B(n1662), .A(n1711), .Z(n1184) );
  CAN2XL U2096 ( .A(n1621), .B(n207), .Z(n1648) );
  COND1X2 U2097 ( .A(n280), .B(n292), .C(n281), .Z(n279) );
  CANR1X2 U2098 ( .A(n312), .B(n293), .C(n294), .Z(n292) );
  COND2XL U2099 ( .A(n77), .B(n1201), .C(n1200), .D(n74), .Z(n922) );
  COND2XL U2100 ( .A(n77), .B(n1202), .C(n1201), .D(n74), .Z(n923) );
  COND2XL U2101 ( .A(n77), .B(n1209), .C(n1208), .D(n74), .Z(n930) );
  COND2XL U2102 ( .A(n77), .B(n1215), .C(n1214), .D(n74), .Z(n936) );
  COND2XL U2103 ( .A(n77), .B(n1208), .C(n1207), .D(n74), .Z(n929) );
  CNR2IXL U2104 ( .B(n1662), .A(n74), .Z(n937) );
  CND2IXL U2105 ( .B(n1661), .A(n1698), .Z(n1235) );
  COND1XL U2106 ( .A(n261), .B(n278), .C(n262), .Z(n260) );
  CENX4 U2107 ( .A(n1688), .B(a[10]), .Z(n50) );
  CND2X4 U2108 ( .A(n1457), .B(n1569), .Z(n18) );
  CND2X4 U2109 ( .A(n1456), .B(n24), .Z(n27) );
  CND2X4 U2110 ( .A(n1455), .B(n33), .Z(n36) );
  CND2X4 U2111 ( .A(n1453), .B(n50), .Z(n53) );
  CIVXL U2112 ( .A(n1670), .Z(n1666) );
  CIVXL U2113 ( .A(n1677), .Z(n1672) );
  CIVXL U2114 ( .A(n1677), .Z(n1673) );
  CIVXL U2115 ( .A(n1677), .Z(n1674) );
  CIVXL U2116 ( .A(n1685), .Z(n1679) );
  CIVXL U2117 ( .A(n1685), .Z(n1680) );
  CIVXL U2118 ( .A(n1684), .Z(n1682) );
  CIVXL U2119 ( .A(n1684), .Z(n1683) );
  CIVXL U2120 ( .A(n1692), .Z(n1686) );
  CIVX1 U2121 ( .A(n93), .Z(n1715) );
  CIVX1 U2122 ( .A(n99), .Z(n1717) );
  CIVX2 U2123 ( .A(n374), .Z(n412) );
  CIVX2 U2124 ( .A(n366), .Z(n410) );
  CIVX2 U2125 ( .A(n358), .Z(n408) );
  CIVX2 U2126 ( .A(n336), .Z(n404) );
  CIVX2 U2127 ( .A(n333), .Z(n403) );
  CIVX2 U2128 ( .A(n322), .Z(n401) );
  CIVX2 U2129 ( .A(n295), .Z(n397) );
  CIVX2 U2130 ( .A(n218), .Z(n387) );
  CIVX2 U2131 ( .A(n380), .Z(n378) );
  CIVX2 U2132 ( .A(n372), .Z(n370) );
  CIVX2 U2133 ( .A(n364), .Z(n362) );
  CIVX2 U2134 ( .A(n356), .Z(n354) );
  CIVX2 U2135 ( .A(n350), .Z(n348) );
  CIVX2 U2136 ( .A(n345), .Z(n343) );
  CIVX2 U2137 ( .A(n339), .Z(n338) );
  CIVX2 U2138 ( .A(n330), .Z(n329) );
  CIVX2 U2139 ( .A(n328), .Z(n326) );
  CIVX2 U2140 ( .A(n327), .Z(n402) );
  CIVX2 U2141 ( .A(n306), .Z(n308) );
  CIVX2 U2142 ( .A(n305), .Z(n399) );
  CIVX2 U2143 ( .A(n303), .Z(n301) );
  CIVX2 U2144 ( .A(n290), .Z(n288) );
  CIVX2 U2145 ( .A(n284), .Z(n395) );
  CIVX2 U2146 ( .A(n279), .Z(n278) );
  CIVX2 U2147 ( .A(n272), .Z(n394) );
  CIVX2 U2148 ( .A(n269), .Z(n393) );
  CIVX2 U2149 ( .A(n261), .Z(n263) );
  CIVX2 U2150 ( .A(n259), .Z(n257) );
  CIVX2 U2151 ( .A(n250), .Z(n248) );
  CIVX2 U2152 ( .A(n249), .Z(n391) );
  CIVX2 U2153 ( .A(n240), .Z(n238) );
  CIVX2 U2154 ( .A(n207), .Z(n205) );
  CIVX2 U2155 ( .A(n104), .Z(n1470) );
  CIVX2 U2156 ( .A(n109), .Z(n1469) );
  CIVX2 U2157 ( .A(n113), .Z(n1468) );
endmodule


module calc_DW_mult_uns_12 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n6, n12, n18, n21, n24, n27, n30, n33, n36, n39, n44, n48, n50, n53,
         n55, n58, n61, n63, n66, n69, n71, n74, n77, n79, n82, n85, n87, n89,
         n91, n93, n95, n97, n99, n100, n102, n104, n105, n107, n109, n110,
         n112, n113, n114, n115, n116, n120, n122, n124, n126, n128, n130,
         n132, n134, n136, n138, n140, n142, n144, n146, n148, n150, n151,
         n152, n153, n154, n155, n156, n157, n169, n170, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n198,
         n199, n205, n207, n208, n210, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n226, n227, n228, n229, n231,
         n234, n235, n236, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n251, n252, n253, n257, n259, n260, n261, n262, n263, n264,
         n268, n270, n271, n272, n273, n275, n278, n279, n280, n281, n283,
         n285, n286, n288, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n301, n303, n304, n305, n306, n308, n311, n312, n313,
         n314, n316, n318, n319, n320, n321, n322, n323, n324, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n343, n345, n346, n348, n350, n351, n352, n354,
         n356, n357, n358, n359, n360, n362, n364, n365, n366, n367, n368,
         n370, n372, n373, n374, n375, n376, n378, n380, n382, n387, n388,
         n389, n390, n394, n397, n399, n401, n402, n403, n404, n408, n410,
         n412, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1455, n1456, n1457, n1468, n1469,
         n1470, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1626,
         n1627, n1628, n1629, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708;
  assign n12 = a[3];
  assign n21 = a[5];
  assign n30 = a[7];
  assign n39 = a[9];
  assign n48 = a[11];
  assign n55 = a[13];
  assign n63 = a[15];
  assign n71 = a[17];
  assign n79 = a[19];
  assign n87 = a[21];
  assign n93 = a[23];
  assign n99 = a[25];
  assign n104 = a[27];
  assign n109 = a[29];
  assign n113 = a[31];
  assign n116 = b[0];
  assign n120 = b[1];
  assign n122 = b[2];
  assign n124 = b[3];
  assign n126 = b[4];
  assign n128 = b[5];
  assign n130 = b[6];
  assign n132 = b[7];
  assign n134 = b[8];
  assign n136 = b[9];
  assign n138 = b[10];
  assign n140 = b[11];
  assign n142 = b[12];
  assign n144 = b[13];
  assign n146 = b[14];
  assign n148 = b[15];
  assign n150 = b[16];
  assign n151 = b[17];
  assign n152 = b[18];
  assign n153 = b[19];
  assign n154 = b[20];
  assign n155 = b[21];
  assign n156 = b[22];
  assign n157 = b[23];

  CNR2X2 U171 ( .A(n513), .B(n538), .Z(n223) );
  CEO3X2 U411 ( .A(n442), .B(n440), .C(n421), .Z(n418) );
  CEO3X2 U412 ( .A(n444), .B(n423), .C(n422), .Z(n419) );
  CEO3X2 U413 ( .A(n425), .B(n424), .C(n446), .Z(n420) );
  CEO3X2 U414 ( .A(n428), .B(n427), .C(n426), .Z(n421) );
  CEO3X2 U415 ( .A(n452), .B(n448), .C(n450), .Z(n422) );
  CEO3X2 U416 ( .A(n429), .B(n456), .C(n454), .Z(n423) );
  CEO3X2 U417 ( .A(n998), .B(n1022), .C(n1106), .Z(n424) );
  CEO3X2 U418 ( .A(n976), .B(n1048), .C(n1076), .Z(n425) );
  CEO3X2 U419 ( .A(n886), .B(n938), .C(n956), .Z(n426) );
  CEO3X2 U420 ( .A(n868), .B(n866), .C(n922), .Z(n427) );
  CEO3X2 U421 ( .A(n872), .B(n896), .C(n908), .Z(n428) );
  CFA1X1 U424 ( .A(n439), .B(n462), .CI(n437), .CO(n432), .S(n433) );
  CFA1X1 U425 ( .A(n441), .B(n464), .CI(n466), .CO(n434), .S(n435) );
  CFA1X1 U426 ( .A(n468), .B(n443), .CI(n445), .CO(n436), .S(n437) );
  CFA1X1 U427 ( .A(n472), .B(n447), .CI(n470), .CO(n438), .S(n439) );
  CFA1X1 U428 ( .A(n474), .B(n449), .CI(n451), .CO(n440), .S(n441) );
  CFA1X1 U429 ( .A(n457), .B(n453), .CI(n455), .CO(n442), .S(n443) );
  CFA1X1 U430 ( .A(n482), .B(n476), .CI(n478), .CO(n444), .S(n445) );
  CFA1X1 U431 ( .A(n999), .B(n480), .CI(n484), .CO(n446), .S(n447) );
  CFA1X1 U432 ( .A(n977), .B(n1107), .CI(n1023), .CO(n448), .S(n449) );
  CFA1X1 U433 ( .A(n957), .B(n1049), .CI(n1077), .CO(n450), .S(n451) );
  CFA1X1 U434 ( .A(n869), .B(n939), .CI(n909), .CO(n452), .S(n453) );
  CFA1X1 U435 ( .A(n887), .B(n923), .CI(n897), .CO(n454), .S(n455) );
  CFA1X1 U437 ( .A(n463), .B(n461), .CI(n488), .CO(n458), .S(n459) );
  CFA1X1 U438 ( .A(n467), .B(n490), .CI(n465), .CO(n460), .S(n461) );
  CFA1X1 U439 ( .A(n469), .B(n492), .CI(n494), .CO(n462), .S(n463) );
  CFA1X1 U440 ( .A(n473), .B(n471), .CI(n496), .CO(n464), .S(n465) );
  CFA1X1 U441 ( .A(n475), .B(n498), .CI(n500), .CO(n466), .S(n467) );
  CFA1X1 U442 ( .A(n481), .B(n477), .CI(n479), .CO(n468), .S(n469) );
  CFA1X1 U443 ( .A(n502), .B(n483), .CI(n504), .CO(n470), .S(n471) );
  CFA1X1 U444 ( .A(n510), .B(n506), .CI(n508), .CO(n472), .S(n473) );
  CFA1X1 U445 ( .A(n1000), .B(n485), .CI(n1024), .CO(n474), .S(n475) );
  CFA1X1 U446 ( .A(n978), .B(n1050), .CI(n1108), .CO(n476), .S(n477) );
  CFA1X1 U447 ( .A(n910), .B(n1078), .CI(n958), .CO(n478), .S(n479) );
  CFA1X1 U448 ( .A(n888), .B(n940), .CI(n898), .CO(n480), .S(n481) );
  CFA1X1 U449 ( .A(n874), .B(n924), .CI(n870), .CO(n482), .S(n483) );
  CHA1X1 U450 ( .A(n851), .B(n880), .CO(n484), .S(n485) );
  CFA1X1 U451 ( .A(n491), .B(n489), .CI(n514), .CO(n486), .S(n487) );
  CFA1X1 U452 ( .A(n495), .B(n516), .CI(n493), .CO(n488), .S(n489) );
  CFA1X1 U453 ( .A(n497), .B(n518), .CI(n520), .CO(n490), .S(n491) );
  CFA1X1 U454 ( .A(n501), .B(n499), .CI(n522), .CO(n492), .S(n493) );
  CFA1X1 U455 ( .A(n503), .B(n524), .CI(n526), .CO(n494), .S(n495) );
  CFA1X1 U456 ( .A(n509), .B(n505), .CI(n507), .CO(n496), .S(n497) );
  CFA1X1 U457 ( .A(n530), .B(n511), .CI(n528), .CO(n498), .S(n499) );
  CFA1X1 U458 ( .A(n536), .B(n534), .CI(n532), .CO(n500), .S(n501) );
  CFA1X1 U459 ( .A(n979), .B(n1025), .CI(n1001), .CO(n502), .S(n503) );
  CFA1X1 U460 ( .A(n959), .B(n1051), .CI(n1109), .CO(n504), .S(n505) );
  CFA1X1 U461 ( .A(n911), .B(n1079), .CI(n925), .CO(n506), .S(n507) );
  CFA1X1 U462 ( .A(n889), .B(n941), .CI(n899), .CO(n508), .S(n509) );
  CFA1X1 U463 ( .A(n871), .B(n875), .CI(n881), .CO(n510), .S(n511) );
  CFA1X1 U464 ( .A(n517), .B(n515), .CI(n540), .CO(n512), .S(n513) );
  CFA1X1 U465 ( .A(n521), .B(n542), .CI(n519), .CO(n514), .S(n515) );
  CFA1X1 U466 ( .A(n546), .B(n544), .CI(n523), .CO(n516), .S(n517) );
  CFA1X1 U467 ( .A(n527), .B(n525), .CI(n548), .CO(n518), .S(n519) );
  CFA1X1 U468 ( .A(n535), .B(n550), .CI(n529), .CO(n520), .S(n521) );
  CFA1X1 U469 ( .A(n552), .B(n531), .CI(n533), .CO(n522), .S(n523) );
  CFA1X1 U470 ( .A(n558), .B(n554), .CI(n556), .CO(n524), .S(n525) );
  CFA1X1 U471 ( .A(n1026), .B(n560), .CI(n537), .CO(n526), .S(n527) );
  CFA1X1 U472 ( .A(n1002), .B(n1080), .CI(n1110), .CO(n528), .S(n529) );
  CFA1X1 U473 ( .A(n926), .B(n1574), .CI(n1629), .CO(n530), .S(n531) );
  CFA1X1 U474 ( .A(n890), .B(n942), .CI(n876), .CO(n532), .S(n533) );
  CFA1X1 U475 ( .A(n900), .B(n960), .CI(n912), .CO(n534), .S(n535) );
  CHA1X1 U476 ( .A(n852), .B(n882), .CO(n536), .S(n537) );
  CFA1X1 U477 ( .A(n543), .B(n541), .CI(n564), .CO(n538), .S(n539) );
  CFA1X1 U478 ( .A(n568), .B(n566), .CI(n545), .CO(n540), .S(n541) );
  CFA1X1 U479 ( .A(n570), .B(n547), .CI(n549), .CO(n542), .S(n543) );
  CFA1X1 U480 ( .A(n574), .B(n551), .CI(n572), .CO(n544), .S(n545) );
  CFA1X1 U481 ( .A(n557), .B(n553), .CI(n555), .CO(n546), .S(n547) );
  CFA1X1 U482 ( .A(n578), .B(n559), .CI(n561), .CO(n548), .S(n549) );
  CFA1X1 U483 ( .A(n582), .B(n576), .CI(n580), .CO(n550), .S(n551) );
  CFA1X1 U486 ( .A(n927), .B(n1081), .CI(n981), .CO(n556), .S(n557) );
  CFA1X1 U488 ( .A(n877), .B(n891), .CI(n883), .CO(n560), .S(n561) );
  CFA1X1 U489 ( .A(n567), .B(n565), .CI(n588), .CO(n562), .S(n563) );
  CFA1X1 U490 ( .A(n592), .B(n590), .CI(n569), .CO(n564), .S(n565) );
  CFA1X1 U491 ( .A(n594), .B(n571), .CI(n573), .CO(n566), .S(n567) );
  CFA1X1 U492 ( .A(n598), .B(n575), .CI(n596), .CO(n568), .S(n569) );
  CFA1X1 U493 ( .A(n581), .B(n577), .CI(n579), .CO(n570), .S(n571) );
  CFA1X1 U494 ( .A(n602), .B(n583), .CI(n600), .CO(n572), .S(n573) );
  CFA1X1 U495 ( .A(n585), .B(n604), .CI(n606), .CO(n574), .S(n575) );
  CFA1X1 U496 ( .A(n962), .B(n1082), .CI(n1112), .CO(n576), .S(n577) );
  CFA1X1 U497 ( .A(n944), .B(n1628), .CI(n1557), .CO(n578), .S(n579) );
  CFA1X1 U498 ( .A(n902), .B(n1004), .CI(n928), .CO(n580), .S(n581) );
  CFA1X1 U499 ( .A(n884), .B(n982), .CI(n914), .CO(n582), .S(n583) );
  CFA1X1 U501 ( .A(n591), .B(n589), .CI(n610), .CO(n586), .S(n587) );
  CFA1X1 U502 ( .A(n614), .B(n593), .CI(n612), .CO(n588), .S(n589) );
  CFA1X1 U503 ( .A(n616), .B(n595), .CI(n597), .CO(n590), .S(n591) );
  CFA1X1 U504 ( .A(n601), .B(n599), .CI(n618), .CO(n592), .S(n593) );
  CFA1X1 U505 ( .A(n605), .B(n620), .CI(n603), .CO(n594), .S(n595) );
  CFA1X1 U506 ( .A(n624), .B(n607), .CI(n622), .CO(n596), .S(n597) );
  CFA1X1 U507 ( .A(n1005), .B(n626), .CI(n628), .CO(n598), .S(n599) );
  CFA1X1 U508 ( .A(n963), .B(n1113), .CI(n1029), .CO(n600), .S(n601) );
  CFA1X1 U509 ( .A(n929), .B(n1083), .CI(n983), .CO(n602), .S(n603) );
  CFA1X1 U511 ( .A(n885), .B(n903), .CI(n893), .CO(n606), .S(n607) );
  CFA1X1 U512 ( .A(n613), .B(n611), .CI(n632), .CO(n608), .S(n609) );
  CFA1X1 U513 ( .A(n617), .B(n634), .CI(n615), .CO(n610), .S(n611) );
  CFA1X1 U515 ( .A(n623), .B(n640), .CI(n621), .CO(n614), .S(n615) );
  CFA1X1 U516 ( .A(n644), .B(n625), .CI(n627), .CO(n616), .S(n617) );
  CFA1X1 U517 ( .A(n648), .B(n642), .CI(n646), .CO(n618), .S(n619) );
  CFA1X1 U518 ( .A(n984), .B(n629), .CI(n1563), .CO(n620), .S(n621) );
  CFA1X1 U519 ( .A(n964), .B(n1056), .CI(n1030), .CO(n622), .S(n623) );
  CFA1X1 U520 ( .A(n916), .B(n1084), .CI(n946), .CO(n624), .S(n625) );
  CFA1X1 U521 ( .A(n894), .B(n1114), .CI(n930), .CO(n626), .S(n627) );
  CFA1X1 U523 ( .A(n635), .B(n633), .CI(n652), .CO(n630), .S(n631) );
  CFA1X1 U524 ( .A(n639), .B(n654), .CI(n637), .CO(n632), .S(n633) );
  CFA1X1 U525 ( .A(n658), .B(n656), .CI(n641), .CO(n634), .S(n635) );
  CFA1X1 U526 ( .A(n645), .B(n660), .CI(n643), .CO(n636), .S(n637) );
  CFA1X1 U527 ( .A(n664), .B(n647), .CI(n649), .CO(n638), .S(n639) );
  CFA1X1 U528 ( .A(n668), .B(n662), .CI(n666), .CO(n640), .S(n641) );
  CFA1X1 U529 ( .A(n965), .B(n1115), .CI(n1007), .CO(n642), .S(n643) );
  CFA1X1 U530 ( .A(n947), .B(n1057), .CI(n1031), .CO(n644), .S(n645) );
  CFA1X1 U531 ( .A(n931), .B(n1085), .CI(n985), .CO(n646), .S(n647) );
  CFA1X1 U532 ( .A(n895), .B(n917), .CI(n905), .CO(n648), .S(n649) );
  CFA1X1 U534 ( .A(n659), .B(n674), .CI(n657), .CO(n652), .S(n653) );
  CFA1X1 U535 ( .A(n678), .B(n676), .CI(n661), .CO(n654), .S(n655) );
  CFA1X1 U536 ( .A(n680), .B(n663), .CI(n665), .CO(n656), .S(n657) );
  CFA1X1 U537 ( .A(n684), .B(n667), .CI(n682), .CO(n658), .S(n659) );
  CFA1X1 U538 ( .A(n986), .B(n686), .CI(n669), .CO(n660), .S(n661) );
  CFA1X1 U539 ( .A(n966), .B(n1058), .CI(n1008), .CO(n662), .S(n663) );
  CFA1X1 U540 ( .A(n948), .B(n1086), .CI(n1032), .CO(n664), .S(n665) );
  CFA1X1 U541 ( .A(n906), .B(n1116), .CI(n932), .CO(n666), .S(n667) );
  CHA1X1 U542 ( .A(n918), .B(n855), .CO(n668), .S(n669) );
  CFA1X1 U543 ( .A(n675), .B(n673), .CI(n690), .CO(n670), .S(n671) );
  CFA1X1 U544 ( .A(n679), .B(n692), .CI(n677), .CO(n672), .S(n673) );
  CFA1X1 U545 ( .A(n681), .B(n694), .CI(n696), .CO(n674), .S(n675) );
  CFA1X1 U546 ( .A(n687), .B(n683), .CI(n685), .CO(n676), .S(n677) );
  CFA1X1 U547 ( .A(n702), .B(n700), .CI(n698), .CO(n678), .S(n679) );
  CFA1X1 U548 ( .A(n987), .B(n704), .CI(n1009), .CO(n680), .S(n681) );
  CFA1X1 U549 ( .A(n967), .B(n1059), .CI(n1117), .CO(n682), .S(n683) );
  CFA1X1 U550 ( .A(n949), .B(n1087), .CI(n1033), .CO(n684), .S(n685) );
  CFA1X1 U551 ( .A(n907), .B(n933), .CI(n919), .CO(n686), .S(n687) );
  CFA1X1 U552 ( .A(n693), .B(n691), .CI(n708), .CO(n688), .S(n689) );
  CFA1X1 U553 ( .A(n697), .B(n710), .CI(n695), .CO(n690), .S(n691) );
  CFA1X1 U554 ( .A(n699), .B(n712), .CI(n714), .CO(n692), .S(n693) );
  CFA1X1 U555 ( .A(n718), .B(n701), .CI(n703), .CO(n694), .S(n695) );
  CFA1X1 U556 ( .A(n705), .B(n716), .CI(n720), .CO(n696), .S(n697) );
  CFA1X1 U557 ( .A(n988), .B(n1010), .CI(n1034), .CO(n698), .S(n699) );
  CFA1X1 U558 ( .A(n968), .B(n1088), .CI(n1118), .CO(n700), .S(n701) );
  CHA1X1 U560 ( .A(n856), .B(n950), .CO(n704), .S(n705) );
  CFA1X1 U561 ( .A(n711), .B(n709), .CI(n724), .CO(n706), .S(n707) );
  CFA1X1 U562 ( .A(n715), .B(n726), .CI(n713), .CO(n708), .S(n709) );
  CFA1X1 U563 ( .A(n717), .B(n728), .CI(n730), .CO(n710), .S(n711) );
  CFA1X1 U564 ( .A(n732), .B(n719), .CI(n721), .CO(n712), .S(n713) );
  CFA1X1 U565 ( .A(n1011), .B(n734), .CI(n736), .CO(n714), .S(n715) );
  CFA1X1 U566 ( .A(n989), .B(n1119), .CI(n1035), .CO(n716), .S(n717) );
  CFA1X1 U567 ( .A(n969), .B(n1089), .CI(n1061), .CO(n718), .S(n719) );
  CFA1X1 U568 ( .A(n921), .B(n951), .CI(n935), .CO(n720), .S(n721) );
  CFA1X1 U569 ( .A(n727), .B(n725), .CI(n740), .CO(n722), .S(n723) );
  CFA1X1 U570 ( .A(n731), .B(n742), .CI(n729), .CO(n724), .S(n725) );
  CFA1X1 U571 ( .A(n735), .B(n744), .CI(n733), .CO(n726), .S(n727) );
  CFA1X1 U572 ( .A(n750), .B(n746), .CI(n748), .CO(n728), .S(n729) );
  CFA1X1 U573 ( .A(n970), .B(n737), .CI(n1120), .CO(n730), .S(n731) );
  CHA1X1 U576 ( .A(n857), .B(n1012), .CO(n736), .S(n737) );
  CFA1X1 U577 ( .A(n743), .B(n741), .CI(n754), .CO(n738), .S(n739) );
  CFA1X1 U578 ( .A(n758), .B(n756), .CI(n745), .CO(n740), .S(n741) );
  CFA1X1 U579 ( .A(n751), .B(n747), .CI(n749), .CO(n742), .S(n743) );
  CFA1X1 U580 ( .A(n764), .B(n762), .CI(n760), .CO(n744), .S(n745) );
  CFA1X1 U581 ( .A(n1013), .B(n1121), .CI(n1037), .CO(n746), .S(n747) );
  CFA1X1 U582 ( .A(n991), .B(n1091), .CI(n1063), .CO(n748), .S(n749) );
  CFA1X1 U583 ( .A(n937), .B(n971), .CI(n953), .CO(n750), .S(n751) );
  CFA1X1 U584 ( .A(n757), .B(n755), .CI(n768), .CO(n752), .S(n753) );
  CFA1X1 U585 ( .A(n772), .B(n759), .CI(n770), .CO(n754), .S(n755) );
  CFA1X1 U586 ( .A(n774), .B(n761), .CI(n763), .CO(n756), .S(n757) );
  CFA1X1 U587 ( .A(n992), .B(n776), .CI(n765), .CO(n758), .S(n759) );
  CFA1X1 U588 ( .A(n972), .B(n1122), .CI(n1014), .CO(n760), .S(n761) );
  CFA1X1 U589 ( .A(n954), .B(n1064), .CI(n1038), .CO(n762), .S(n763) );
  CHA1X1 U590 ( .A(n858), .B(n1092), .CO(n764), .S(n765) );
  CFA1X1 U591 ( .A(n771), .B(n769), .CI(n780), .CO(n766), .S(n767) );
  CFA1X1 U592 ( .A(n775), .B(n782), .CI(n773), .CO(n768), .S(n769) );
  CFA1X1 U593 ( .A(n784), .B(n777), .CI(n786), .CO(n770), .S(n771) );
  CFA1X1 U594 ( .A(n1039), .B(n788), .CI(n1123), .CO(n772), .S(n773) );
  CFA1X1 U595 ( .A(n1015), .B(n1065), .CI(n1093), .CO(n774), .S(n775) );
  CFA1X1 U597 ( .A(n783), .B(n781), .CI(n792), .CO(n778), .S(n779) );
  CFA1X1 U598 ( .A(n787), .B(n794), .CI(n785), .CO(n780), .S(n781) );
  CFA1X1 U599 ( .A(n789), .B(n796), .CI(n798), .CO(n782), .S(n783) );
  CFA1X1 U600 ( .A(n994), .B(n1040), .CI(n1016), .CO(n784), .S(n785) );
  CFA1X1 U601 ( .A(n974), .B(n1066), .CI(n1124), .CO(n786), .S(n787) );
  CHA1X1 U602 ( .A(n859), .B(n1094), .CO(n788), .S(n789) );
  CFA1X1 U603 ( .A(n802), .B(n793), .CI(n795), .CO(n790), .S(n791) );
  CFA1X1 U604 ( .A(n799), .B(n804), .CI(n797), .CO(n792), .S(n793) );
  CFA1X1 U605 ( .A(n1125), .B(n806), .CI(n808), .CO(n794), .S(n795) );
  CFA1X1 U607 ( .A(n975), .B(n1017), .CI(n995), .CO(n798), .S(n799) );
  CFA1X1 U608 ( .A(n805), .B(n803), .CI(n812), .CO(n800), .S(n801) );
  CFA1X1 U609 ( .A(n816), .B(n807), .CI(n814), .CO(n802), .S(n803) );
  CFA1X1 U610 ( .A(n1018), .B(n809), .CI(n1042), .CO(n804), .S(n805) );
  CFA1X1 U611 ( .A(n996), .B(n1068), .CI(n1126), .CO(n806), .S(n807) );
  CHA1X1 U612 ( .A(n860), .B(n1096), .CO(n808), .S(n809) );
  CFA1X1 U613 ( .A(n815), .B(n813), .CI(n820), .CO(n810), .S(n811) );
  CFA1X1 U614 ( .A(n824), .B(n817), .CI(n822), .CO(n812), .S(n813) );
  CFA1X1 U615 ( .A(n1127), .B(n1097), .CI(n1069), .CO(n814), .S(n815) );
  CFA1X1 U616 ( .A(n997), .B(n1043), .CI(n1019), .CO(n816), .S(n817) );
  CFA1X1 U617 ( .A(n828), .B(n821), .CI(n823), .CO(n818), .S(n819) );
  CFA1X1 U618 ( .A(n1044), .B(n830), .CI(n825), .CO(n820), .S(n821) );
  CFA1X1 U619 ( .A(n1020), .B(n1070), .CI(n1128), .CO(n822), .S(n823) );
  CHA1X1 U620 ( .A(n861), .B(n1098), .CO(n824), .S(n825) );
  CFA1X1 U621 ( .A(n834), .B(n829), .CI(n831), .CO(n826), .S(n827) );
  CFA1X1 U622 ( .A(n1099), .B(n836), .CI(n1071), .CO(n828), .S(n829) );
  CFA1X1 U623 ( .A(n1021), .B(n1129), .CI(n1045), .CO(n830), .S(n831) );
  CFA1X1 U624 ( .A(n837), .B(n835), .CI(n840), .CO(n832), .S(n833) );
  CFA1X1 U625 ( .A(n1046), .B(n1072), .CI(n1130), .CO(n834), .S(n835) );
  CHA1X1 U626 ( .A(n862), .B(n1100), .CO(n836), .S(n837) );
  CFA1X1 U627 ( .A(n1073), .B(n841), .CI(n844), .CO(n838), .S(n839) );
  CFA1X1 U628 ( .A(n1047), .B(n1101), .CI(n1131), .CO(n840), .S(n841) );
  CFA1X1 U629 ( .A(n1102), .B(n845), .CI(n1074), .CO(n842), .S(n843) );
  CHA1X1 U630 ( .A(n1132), .B(n863), .CO(n844), .S(n845) );
  CFA1X1 U631 ( .A(n1075), .B(n1103), .CI(n1133), .CO(n846), .S(n847) );
  CHA1X1 U632 ( .A(n1134), .B(n1104), .CO(n848), .S(n849) );
  COND2X1 U633 ( .A(n115), .B(n1468), .C(n114), .D(n1139), .Z(n850) );
  COND2X1 U634 ( .A(n1137), .B(n114), .C(n115), .D(n1138), .Z(n866) );
  CND2IX1 U638 ( .B(n1706), .A(n113), .Z(n1139) );
  COND2X1 U639 ( .A(n112), .B(n1469), .C(n110), .D(n1144), .Z(n851) );
  COND2X1 U640 ( .A(n1140), .B(n110), .C(n1141), .D(n112), .Z(n868) );
  COND2X1 U641 ( .A(n1142), .B(n112), .C(n110), .D(n1141), .Z(n869) );
  COND2X1 U642 ( .A(n1142), .B(n110), .C(n112), .D(n1143), .Z(n870) );
  CND2IX1 U648 ( .B(n1706), .A(n109), .Z(n1144) );
  COND2X1 U649 ( .A(n107), .B(n1470), .C(n105), .D(n1151), .Z(n852) );
  COND2X1 U650 ( .A(n1145), .B(n105), .C(n1146), .D(n107), .Z(n872) );
  COND2X1 U652 ( .A(n1147), .B(n105), .C(n1148), .D(n107), .Z(n874) );
  COND2X1 U653 ( .A(n1149), .B(n107), .C(n105), .D(n1148), .Z(n875) );
  COND2X1 U654 ( .A(n1149), .B(n105), .C(n107), .D(n1150), .Z(n876) );
  CND2IX1 U662 ( .B(n1706), .A(n104), .Z(n1151) );
  CND2IX1 U680 ( .B(n1706), .A(n1703), .Z(n1160) );
  COND2X1 U683 ( .A(n97), .B(n1163), .C(n1162), .D(n95), .Z(n887) );
  COND2X1 U684 ( .A(n97), .B(n1164), .C(n95), .D(n1163), .Z(n888) );
  COND2X1 U685 ( .A(n1165), .B(n97), .C(n1164), .D(n95), .Z(n889) );
  COND2X1 U686 ( .A(n1165), .B(n95), .C(n1166), .D(n97), .Z(n890) );
  COND2X1 U689 ( .A(n1169), .B(n97), .C(n1168), .D(n95), .Z(n893) );
  COND2X1 U690 ( .A(n1170), .B(n97), .C(n95), .D(n1169), .Z(n894) );
  COND2X1 U703 ( .A(n91), .B(n1700), .C(n1184), .D(n89), .Z(n855) );
  COND2X1 U704 ( .A(n91), .B(n1173), .C(n89), .D(n1172), .Z(n896) );
  COND2X1 U705 ( .A(n91), .B(n1174), .C(n1173), .D(n89), .Z(n897) );
  COND2X1 U706 ( .A(n91), .B(n1175), .C(n89), .D(n1174), .Z(n898) );
  COND2X1 U707 ( .A(n91), .B(n1176), .C(n1175), .D(n89), .Z(n899) );
  COND2X1 U708 ( .A(n91), .B(n1177), .C(n89), .D(n1176), .Z(n900) );
  COND2X1 U710 ( .A(n91), .B(n1179), .C(n89), .D(n1178), .Z(n902) );
  COND2X1 U712 ( .A(n91), .B(n1181), .C(n89), .D(n1180), .Z(n904) );
  COND2X1 U713 ( .A(n91), .B(n1182), .C(n1181), .D(n89), .Z(n905) );
  COND2X1 U714 ( .A(n91), .B(n1183), .C(n89), .D(n1182), .Z(n906) );
  CND2IX1 U728 ( .B(n1706), .A(n1698), .Z(n1184) );
  COND2X1 U736 ( .A(n1633), .B(n1192), .C(n82), .D(n1191), .Z(n914) );
  CND2IX1 U758 ( .B(n1706), .A(n1694), .Z(n1199) );
  COND2X1 U761 ( .A(n77), .B(n1202), .C(n1201), .D(n74), .Z(n923) );
  COND2X1 U762 ( .A(n77), .B(n1203), .C(n1202), .D(n74), .Z(n924) );
  COND2X1 U763 ( .A(n77), .B(n1204), .C(n1203), .D(n74), .Z(n925) );
  COND2X1 U764 ( .A(n77), .B(n1205), .C(n1204), .D(n74), .Z(n926) );
  COND2X1 U765 ( .A(n77), .B(n1206), .C(n1205), .D(n74), .Z(n927) );
  COND2X1 U766 ( .A(n77), .B(n1207), .C(n1206), .D(n74), .Z(n928) );
  COND2X1 U767 ( .A(n77), .B(n1208), .C(n1207), .D(n74), .Z(n929) );
  COND2X1 U768 ( .A(n77), .B(n1209), .C(n74), .D(n1208), .Z(n930) );
  COND2X1 U769 ( .A(n77), .B(n1210), .C(n1209), .D(n74), .Z(n931) );
  COND2X1 U770 ( .A(n77), .B(n1211), .C(n74), .D(n1210), .Z(n932) );
  COND2X1 U773 ( .A(n77), .B(n1214), .C(n1213), .D(n74), .Z(n935) );
  COND2X1 U774 ( .A(n77), .B(n1215), .C(n74), .D(n1214), .Z(n936) );
  COND2X1 U800 ( .A(n69), .B(n1224), .C(n1223), .D(n66), .Z(n944) );
  COND2X1 U801 ( .A(n69), .B(n1225), .C(n1224), .D(n66), .Z(n945) );
  COND2X1 U803 ( .A(n69), .B(n1227), .C(n1226), .D(n66), .Z(n947) );
  COND2X1 U804 ( .A(n69), .B(n1228), .C(n1227), .D(n66), .Z(n948) );
  COND2X1 U805 ( .A(n69), .B(n1229), .C(n1228), .D(n66), .Z(n949) );
  COND2X1 U807 ( .A(n69), .B(n1231), .C(n1230), .D(n66), .Z(n951) );
  COND2X1 U809 ( .A(n69), .B(n1233), .C(n1232), .D(n66), .Z(n953) );
  COND2X1 U810 ( .A(n69), .B(n1234), .C(n66), .D(n1233), .Z(n954) );
  COND2X1 U831 ( .A(n61), .B(n1560), .C(n1256), .D(n58), .Z(n859) );
  COND2X1 U832 ( .A(n61), .B(n1237), .C(n1236), .D(n58), .Z(n956) );
  COND2X1 U833 ( .A(n61), .B(n1238), .C(n1237), .D(n58), .Z(n957) );
  COND2X1 U834 ( .A(n61), .B(n1239), .C(n1238), .D(n58), .Z(n958) );
  COND2X1 U835 ( .A(n61), .B(n1240), .C(n1239), .D(n58), .Z(n959) );
  COND2X1 U836 ( .A(n61), .B(n1241), .C(n1240), .D(n58), .Z(n960) );
  COND2X1 U837 ( .A(n61), .B(n1242), .C(n1241), .D(n58), .Z(n961) );
  COND2X1 U838 ( .A(n61), .B(n1243), .C(n1242), .D(n58), .Z(n962) );
  COND2X1 U839 ( .A(n61), .B(n1244), .C(n1243), .D(n58), .Z(n963) );
  COND2X1 U840 ( .A(n61), .B(n1245), .C(n1244), .D(n58), .Z(n964) );
  COND2X1 U841 ( .A(n61), .B(n1246), .C(n1245), .D(n58), .Z(n965) );
  COND2X1 U842 ( .A(n61), .B(n1247), .C(n1246), .D(n58), .Z(n966) );
  COND2X1 U843 ( .A(n61), .B(n1248), .C(n1247), .D(n58), .Z(n967) );
  COND2X1 U844 ( .A(n61), .B(n1249), .C(n1248), .D(n58), .Z(n968) );
  COND2X1 U845 ( .A(n61), .B(n1250), .C(n1249), .D(n58), .Z(n969) );
  COND2X1 U846 ( .A(n61), .B(n1251), .C(n58), .D(n1250), .Z(n970) );
  COND2X1 U847 ( .A(n61), .B(n1252), .C(n1251), .D(n58), .Z(n971) );
  COND2X1 U848 ( .A(n61), .B(n1253), .C(n58), .D(n1252), .Z(n972) );
  COND2X1 U849 ( .A(n61), .B(n1254), .C(n1253), .D(n58), .Z(n973) );
  COND2X1 U850 ( .A(n61), .B(n1255), .C(n58), .D(n1254), .Z(n974) );
  CND2IX1 U872 ( .B(n1706), .A(n1684), .Z(n1256) );
  COND2X1 U880 ( .A(n53), .B(n1264), .C(n1263), .D(n50), .Z(n982) );
  COND2X1 U883 ( .A(n53), .B(n1267), .C(n1266), .D(n50), .Z(n985) );
  COND2X1 U889 ( .A(n53), .B(n1273), .C(n1272), .D(n50), .Z(n991) );
  COND2X1 U926 ( .A(n44), .B(n1287), .C(n1286), .D(n1559), .Z(n1004) );
  COND2X1 U929 ( .A(n44), .B(n1290), .C(n1289), .D(n1559), .Z(n1007) );
  COND2X1 U930 ( .A(n44), .B(n1291), .C(n1290), .D(n1559), .Z(n1008) );
  COND2X1 U935 ( .A(n44), .B(n1296), .C(n1295), .D(n1559), .Z(n1013) );
  COND2X1 U936 ( .A(n44), .B(n1297), .C(n1296), .D(n1559), .Z(n1014) );
  COND2X1 U941 ( .A(n44), .B(n1302), .C(n1301), .D(n1559), .Z(n1019) );
  COND2X1 U977 ( .A(n36), .B(n1313), .C(n1312), .D(n33), .Z(n1029) );
  COND2X1 U979 ( .A(n36), .B(n1315), .C(n1314), .D(n33), .Z(n1031) );
  COND2X1 U980 ( .A(n36), .B(n1316), .C(n1315), .D(n33), .Z(n1032) );
  COND2X1 U981 ( .A(n36), .B(n1317), .C(n1316), .D(n33), .Z(n1033) );
  COND2X1 U985 ( .A(n36), .B(n1321), .C(n1320), .D(n33), .Z(n1037) );
  COND2X1 U986 ( .A(n36), .B(n1322), .C(n1321), .D(n33), .Z(n1038) );
  CND2IX1 U1022 ( .B(n1706), .A(n1669), .Z(n1331) );
  COND2X1 U1023 ( .A(n27), .B(n1665), .C(n1360), .D(n24), .Z(n863) );
  COND2X1 U1024 ( .A(n27), .B(n1333), .C(n24), .D(n1332), .Z(n1048) );
  COND2X1 U1025 ( .A(n27), .B(n1334), .C(n24), .D(n1333), .Z(n1049) );
  COND2X1 U1026 ( .A(n27), .B(n1335), .C(n24), .D(n1334), .Z(n1050) );
  COND2X1 U1027 ( .A(n27), .B(n1336), .C(n24), .D(n1335), .Z(n1051) );
  COND2X1 U1029 ( .A(n27), .B(n1338), .C(n24), .D(n1337), .Z(n1053) );
  COND2X1 U1031 ( .A(n27), .B(n1340), .C(n24), .D(n1339), .Z(n1055) );
  COND2X1 U1033 ( .A(n27), .B(n1342), .C(n24), .D(n1341), .Z(n1057) );
  COND2X1 U1034 ( .A(n27), .B(n1343), .C(n24), .D(n1342), .Z(n1058) );
  COND2X1 U1035 ( .A(n27), .B(n1344), .C(n24), .D(n1343), .Z(n1059) );
  COND2X1 U1036 ( .A(n27), .B(n1345), .C(n24), .D(n1344), .Z(n1060) );
  COND2X1 U1037 ( .A(n27), .B(n1346), .C(n24), .D(n1345), .Z(n1061) );
  COND2X1 U1038 ( .A(n27), .B(n1347), .C(n24), .D(n1346), .Z(n1062) );
  COND2X1 U1039 ( .A(n27), .B(n1348), .C(n24), .D(n1347), .Z(n1063) );
  COND2X1 U1040 ( .A(n27), .B(n1349), .C(n24), .D(n1348), .Z(n1064) );
  COND2X1 U1041 ( .A(n27), .B(n1350), .C(n24), .D(n1349), .Z(n1065) );
  COND2X1 U1042 ( .A(n27), .B(n1351), .C(n24), .D(n1350), .Z(n1066) );
  COND2X1 U1043 ( .A(n27), .B(n1352), .C(n24), .D(n1351), .Z(n1067) );
  COND2X1 U1044 ( .A(n27), .B(n1353), .C(n24), .D(n1352), .Z(n1068) );
  COND2X1 U1045 ( .A(n27), .B(n1354), .C(n24), .D(n1353), .Z(n1069) );
  COND2X1 U1046 ( .A(n27), .B(n1355), .C(n24), .D(n1354), .Z(n1070) );
  COND2X1 U1047 ( .A(n27), .B(n1356), .C(n24), .D(n1355), .Z(n1071) );
  COND2X1 U1048 ( .A(n27), .B(n1357), .C(n24), .D(n1356), .Z(n1072) );
  COND2X1 U1049 ( .A(n27), .B(n1358), .C(n24), .D(n1357), .Z(n1073) );
  COND2X1 U1050 ( .A(n27), .B(n1359), .C(n24), .D(n1358), .Z(n1074) );
  COND2X1 U1084 ( .A(n18), .B(n1364), .C(n1626), .D(n1363), .Z(n1078) );
  COND2X1 U1085 ( .A(n18), .B(n1365), .C(n1626), .D(n1364), .Z(n1079) );
  COND2X1 U1086 ( .A(n18), .B(n1366), .C(n1626), .D(n1365), .Z(n1080) );
  COND2X1 U1087 ( .A(n18), .B(n1367), .C(n1626), .D(n1366), .Z(n1081) );
  COND2X1 U1088 ( .A(n18), .B(n1368), .C(n1626), .D(n1367), .Z(n1082) );
  COND2X1 U1089 ( .A(n18), .B(n1369), .C(n1626), .D(n1368), .Z(n1083) );
  COND2X1 U1090 ( .A(n18), .B(n1370), .C(n1626), .D(n1369), .Z(n1084) );
  COND2X1 U1091 ( .A(n18), .B(n1371), .C(n1626), .D(n1370), .Z(n1085) );
  COND2X1 U1092 ( .A(n18), .B(n1372), .C(n1626), .D(n1371), .Z(n1086) );
  COND2X1 U1093 ( .A(n18), .B(n1373), .C(n1626), .D(n1372), .Z(n1087) );
  COND2X1 U1094 ( .A(n18), .B(n1374), .C(n1626), .D(n1373), .Z(n1088) );
  COND2X1 U1095 ( .A(n18), .B(n1375), .C(n1626), .D(n1374), .Z(n1089) );
  COND2X1 U1096 ( .A(n18), .B(n1376), .C(n1626), .D(n1375), .Z(n1090) );
  COND2X1 U1097 ( .A(n18), .B(n1377), .C(n1626), .D(n1376), .Z(n1091) );
  COND2X1 U1099 ( .A(n18), .B(n1379), .C(n1626), .D(n1378), .Z(n1093) );
  COND2X1 U1100 ( .A(n18), .B(n1380), .C(n1626), .D(n1379), .Z(n1094) );
  COND2X1 U1101 ( .A(n18), .B(n1381), .C(n1626), .D(n1380), .Z(n1095) );
  COND2X1 U1103 ( .A(n18), .B(n1383), .C(n1626), .D(n1382), .Z(n1097) );
  COND2X1 U1104 ( .A(n18), .B(n1384), .C(n1626), .D(n1383), .Z(n1098) );
  COND2X1 U1106 ( .A(n18), .B(n1386), .C(n1626), .D(n1385), .Z(n1100) );
  COND2X1 U1109 ( .A(n18), .B(n1389), .C(n1626), .D(n1388), .Z(n1103) );
  COND2X1 U1110 ( .A(n18), .B(n1390), .C(n1626), .D(n1389), .Z(n1104) );
  CEOX2 U1241 ( .A(a[24]), .B(n1703), .Z(n1446) );
  CEOX2 U1268 ( .A(a[6]), .B(n1670), .Z(n1455) );
  CNR2X2 U1281 ( .A(n6), .B(n1392), .Z(n1106) );
  CNR2X2 U1282 ( .A(n6), .B(n1395), .Z(n1109) );
  CNR2X2 U1283 ( .A(n6), .B(n1397), .Z(n1111) );
  CNR2X2 U1284 ( .A(n6), .B(n1399), .Z(n1113) );
  CNR2X2 U1285 ( .A(n6), .B(n1400), .Z(n1114) );
  CNR2X2 U1286 ( .A(n6), .B(n1413), .Z(n1127) );
  CNR2X2 U1287 ( .A(n6), .B(n1414), .Z(n1128) );
  CNR2X2 U1288 ( .A(n6), .B(n1415), .Z(n1129) );
  CNR2X2 U1289 ( .A(n6), .B(n1420), .Z(n1134) );
  CNR2X2 U1290 ( .A(n6), .B(n1421), .Z(n1135) );
  CNR2X2 U1291 ( .A(n6), .B(n1422), .Z(n1136) );
  CNR2X2 U1292 ( .A(n6), .B(n1412), .Z(n1126) );
  CNR2X2 U1293 ( .A(n6), .B(n1411), .Z(n1125) );
  CNR2X2 U1294 ( .A(n6), .B(n1410), .Z(n1124) );
  CNR2X2 U1295 ( .A(n6), .B(n1408), .Z(n1122) );
  CNR2X2 U1296 ( .A(n6), .B(n1405), .Z(n1119) );
  CNR2X2 U1297 ( .A(n6), .B(n1402), .Z(n1116) );
  CNR2X2 U1298 ( .A(n6), .B(n1396), .Z(n1110) );
  CNR2X2 U1299 ( .A(n6), .B(n1417), .Z(n1131) );
  CNR2X2 U1300 ( .A(n6), .B(n1418), .Z(n1132) );
  CNR2X2 U1301 ( .A(n6), .B(n1419), .Z(n1133) );
  CNR2X2 U1302 ( .A(n6), .B(n1407), .Z(n1121) );
  CNR2X2 U1303 ( .A(n6), .B(n1404), .Z(n1118) );
  CNR2X2 U1304 ( .A(n6), .B(n1403), .Z(n1117) );
  CNR2X2 U1305 ( .A(n6), .B(n1401), .Z(n1115) );
  CNR2X2 U1306 ( .A(n6), .B(n1393), .Z(n1107) );
  CNR2X2 U1307 ( .A(n6), .B(n1394), .Z(n1108) );
  CNR2X2 U1308 ( .A(n6), .B(n1416), .Z(n1130) );
  CNR2X2 U1309 ( .A(n6), .B(n1406), .Z(n1120) );
  CNR2X2 U1310 ( .A(n6), .B(n1409), .Z(n1123) );
  CNR2X2 U1311 ( .A(n6), .B(n1398), .Z(n1112) );
  CIVX2 U1312 ( .A(b[31]), .Z(n1392) );
  CIVX2 U1313 ( .A(n1651), .Z(n1414) );
  CIVX2 U1314 ( .A(n1652), .Z(n1413) );
  CIVX2 U1315 ( .A(n142), .Z(n1411) );
  CIVX2 U1316 ( .A(n1653), .Z(n1412) );
  CIVX2 U1317 ( .A(n1648), .Z(n1417) );
  CIVX2 U1318 ( .A(n1647), .Z(n1418) );
  CIVX2 U1319 ( .A(n1644), .Z(n1421) );
  CENXL U1320 ( .A(1'b0), .B(n148), .Z(n1408) );
  CENXL U1321 ( .A(1'b0), .B(n1646), .Z(n1419) );
  CIVX2 U1322 ( .A(n1650), .Z(n1415) );
  CIVX2 U1323 ( .A(b[30]), .Z(n1393) );
  CIVX2 U1324 ( .A(b[28]), .Z(n1395) );
  CIVX2 U1325 ( .A(b[27]), .Z(n1396) );
  CIVX2 U1326 ( .A(b[26]), .Z(n1397) );
  CIVX2 U1327 ( .A(b[24]), .Z(n1399) );
  CIVX2 U1328 ( .A(n156), .Z(n1401) );
  CIVX2 U1329 ( .A(n154), .Z(n1403) );
  CIVX2 U1330 ( .A(n155), .Z(n1402) );
  CENXL U1331 ( .A(1'b0), .B(b[25]), .Z(n1398) );
  CENXL U1332 ( .A(1'b0), .B(b[29]), .Z(n1394) );
  CIVX2 U1333 ( .A(n157), .Z(n1400) );
  CIVX2 U1334 ( .A(n153), .Z(n1404) );
  CENXL U1335 ( .A(1'b0), .B(n1649), .Z(n1416) );
  CIVX2 U1336 ( .A(n150), .Z(n1407) );
  CIVX2 U1337 ( .A(n146), .Z(n1409) );
  CIVX2 U1338 ( .A(n1707), .Z(n1422) );
  CIVX2 U1339 ( .A(n1654), .Z(n1410) );
  CIVX2 U1340 ( .A(n151), .Z(n1406) );
  CIVX2 U1341 ( .A(n1645), .Z(n1420) );
  CENXL U1342 ( .A(1'b0), .B(n152), .Z(n1405) );
  CIVX2 U1343 ( .A(n1136), .Z(n382) );
  CIVX2 U1344 ( .A(n382), .Z(product[1]) );
  CIVX2 U1345 ( .A(n195), .Z(product[2]) );
  CIVX2 U1346 ( .A(n378), .Z(n376) );
  CIVX2 U1347 ( .A(n1665), .Z(n1662) );
  CIVX3 U1348 ( .A(n1704), .Z(n1703) );
  CND2X2 U1349 ( .A(n1445), .B(n105), .Z(n107) );
  CENX1 U1350 ( .A(n1705), .B(n104), .Z(n1150) );
  CENXL U1351 ( .A(n1707), .B(n1678), .Z(n1302) );
  CND2X4 U1352 ( .A(n95), .B(n1447), .Z(n97) );
  COND2X1 U1353 ( .A(n36), .B(n1320), .C(n1319), .D(n33), .Z(n1036) );
  CND2X4 U1354 ( .A(n1455), .B(n33), .Z(n36) );
  CIVX3 U1355 ( .A(n21), .Z(n1665) );
  CIVX2 U1356 ( .A(n1665), .Z(n1664) );
  CIVX4 U1357 ( .A(n1665), .Z(n1663) );
  CENXL U1358 ( .A(n1677), .B(n1654), .Z(n1290) );
  CNIVX1 U1359 ( .A(n1028), .Z(n1557) );
  CENXL U1360 ( .A(n1681), .B(n153), .Z(n1259) );
  CENXL U1361 ( .A(n1647), .B(n1681), .Z(n1273) );
  CENXL U1362 ( .A(n1645), .B(n1681), .Z(n1275) );
  CENXL U1363 ( .A(n1707), .B(n1681), .Z(n1277) );
  CENXL U1364 ( .A(n1681), .B(n1652), .Z(n1268) );
  CENXL U1365 ( .A(n1684), .B(n152), .Z(n1237) );
  CENXL U1366 ( .A(n1681), .B(n152), .Z(n1260) );
  CENXL U1367 ( .A(n1664), .B(n152), .Z(n1341) );
  CENXL U1368 ( .A(n1701), .B(n1650), .Z(n1162) );
  CENXL U1369 ( .A(n1698), .B(n1650), .Z(n1175) );
  CENXL U1370 ( .A(n1658), .B(n1650), .Z(n1382) );
  CENXL U1371 ( .A(n1675), .B(n1650), .Z(n1295) );
  CENXL U1372 ( .A(n1663), .B(n1650), .Z(n1351) );
  CENXL U1373 ( .A(n1681), .B(n1650), .Z(n1270) );
  CENXL U1374 ( .A(n1646), .B(n104), .Z(n1146) );
  CENXL U1375 ( .A(n1674), .B(n1646), .Z(n1299) );
  CENXL U1376 ( .A(n1646), .B(n1703), .Z(n1155) );
  CENXL U1377 ( .A(n1681), .B(n1646), .Z(n1274) );
  CENXL U1378 ( .A(n1699), .B(n1646), .Z(n1179) );
  CENXL U1379 ( .A(n1693), .B(n1646), .Z(n1194) );
  CENXL U1380 ( .A(n1705), .B(n113), .Z(n1138) );
  CENXL U1381 ( .A(n1705), .B(n109), .Z(n1143) );
  CENXL U1382 ( .A(n1705), .B(n1674), .Z(n1303) );
  CENXL U1383 ( .A(n1705), .B(n1681), .Z(n1278) );
  CENXL U1384 ( .A(n1705), .B(n1690), .Z(n1215) );
  CENXL U1385 ( .A(n1705), .B(n1686), .Z(n1234) );
  CENXL U1386 ( .A(n1705), .B(n1699), .Z(n1183) );
  CENXL U1387 ( .A(n1705), .B(n1703), .Z(n1159) );
  CENX1 U1388 ( .A(n1705), .B(n1701), .Z(n1170) );
  CENXL U1389 ( .A(n1649), .B(n1703), .Z(n1152) );
  CENXL U1390 ( .A(n1657), .B(n1649), .Z(n1383) );
  CENXL U1391 ( .A(n1649), .B(n1701), .Z(n1163) );
  CENXL U1392 ( .A(n1666), .B(n1649), .Z(n1323) );
  CENXL U1393 ( .A(n1649), .B(n1699), .Z(n1176) );
  CENXL U1394 ( .A(n1664), .B(n1649), .Z(n1352) );
  CENXL U1395 ( .A(n1649), .B(n1686), .Z(n1227) );
  CENXL U1396 ( .A(n1681), .B(n1649), .Z(n1271) );
  CENXL U1397 ( .A(n1649), .B(n1689), .Z(n1208) );
  CENX1 U1398 ( .A(n1649), .B(n1694), .Z(n1191) );
  COND1XL U1399 ( .A(n376), .B(n374), .C(n375), .Z(n373) );
  CNIVX2 U1400 ( .A(n128), .Z(n1647) );
  CENX1 U1401 ( .A(n1659), .B(n150), .Z(n1374) );
  CENX1 U1402 ( .A(n1645), .B(n1699), .Z(n1180) );
  CENX1 U1403 ( .A(n1681), .B(n146), .Z(n1264) );
  CENX1 U1404 ( .A(n1645), .B(n1701), .Z(n1167) );
  CENX1 U1405 ( .A(n1688), .B(n1650), .Z(n1207) );
  CENX1 U1406 ( .A(n1668), .B(n152), .Z(n1312) );
  CENX1 U1407 ( .A(n1646), .B(n1701), .Z(n1166) );
  CENX1 U1408 ( .A(n1669), .B(n153), .Z(n1311) );
  CENX1 U1409 ( .A(n1681), .B(n150), .Z(n1262) );
  CENX1 U1410 ( .A(n1681), .B(n148), .Z(n1263) );
  CENX1 U1411 ( .A(n1693), .B(n1650), .Z(n1190) );
  CENX1 U1412 ( .A(n1677), .B(n150), .Z(n1287) );
  CENX1 U1413 ( .A(n1707), .B(n1701), .Z(n1169) );
  CENX1 U1414 ( .A(n1681), .B(n1654), .Z(n1265) );
  CENX1 U1415 ( .A(n1645), .B(n1686), .Z(n1231) );
  CENX1 U1416 ( .A(n1664), .B(n1654), .Z(n1346) );
  CENX1 U1417 ( .A(n1707), .B(n1689), .Z(n1214) );
  CENX1 U1418 ( .A(n1681), .B(n1648), .Z(n1272) );
  CENX1 U1419 ( .A(n1645), .B(n1703), .Z(n1156) );
  CENX1 U1420 ( .A(n1686), .B(n1654), .Z(n1221) );
  CENX1 U1421 ( .A(n1647), .B(n1701), .Z(n1165) );
  CENX1 U1422 ( .A(n1673), .B(n153), .Z(n1284) );
  CENX1 U1423 ( .A(n1664), .B(b[24]), .Z(n1335) );
  CENX1 U1424 ( .A(n1701), .B(n1648), .Z(n1164) );
  CENX1 U1425 ( .A(n1658), .B(n153), .Z(n1371) );
  CENX1 U1426 ( .A(n1681), .B(n1653), .Z(n1267) );
  CENX1 U1427 ( .A(n1681), .B(n142), .Z(n1266) );
  COR2X1 U1428 ( .A(n1578), .B(n1579), .Z(n918) );
  CND3XL U1429 ( .A(n1637), .B(n1638), .C(n1639), .Z(n702) );
  CENX1 U1430 ( .A(n1645), .B(n1678), .Z(n1300) );
  CENX1 U1431 ( .A(n1645), .B(n104), .Z(n1147) );
  CENX1 U1432 ( .A(n1703), .B(a[26]), .Z(n105) );
  CEOX1 U1433 ( .A(a[26]), .B(n104), .Z(n1445) );
  CENX1 U1434 ( .A(n1657), .B(b[27]), .Z(n1363) );
  CENX1 U1435 ( .A(n1663), .B(b[26]), .Z(n1333) );
  CENX1 U1436 ( .A(n1645), .B(n1670), .Z(n1327) );
  CNIVX2 U1437 ( .A(n1601), .Z(n1559) );
  CIVX4 U1438 ( .A(n1623), .Z(n33) );
  CEOX2 U1439 ( .A(n1663), .B(a[6]), .Z(n1623) );
  CND2X1 U1440 ( .A(n1592), .B(n1593), .Z(n879) );
  CENX1 U1441 ( .A(n1645), .B(n109), .Z(n1140) );
  CENX1 U1442 ( .A(n1707), .B(n1659), .Z(n1389) );
  CENX1 U1443 ( .A(n1657), .B(n1645), .Z(n1387) );
  CIVX4 U1444 ( .A(a[2]), .Z(n1626) );
  CEOX1 U1445 ( .A(a[4]), .B(n1663), .Z(n1456) );
  CEOX1 U1446 ( .A(n1594), .B(n433), .Z(n431) );
  CEOX1 U1447 ( .A(n435), .B(n460), .Z(n1594) );
  CANR1X1 U1448 ( .A(n288), .B(n1611), .C(n283), .Z(n281) );
  CNR2X1 U1449 ( .A(n707), .B(n722), .Z(n295) );
  CANR1X1 U1450 ( .A(n308), .B(n1612), .C(n301), .Z(n299) );
  CNIVX2 U1451 ( .A(n116), .Z(n1706) );
  CND2X1 U1452 ( .A(n459), .B(n486), .Z(n212) );
  CND3XL U1453 ( .A(n1595), .B(n1596), .C(n1597), .Z(n430) );
  CND2X1 U1454 ( .A(n431), .B(n458), .Z(n207) );
  CANR1XL U1455 ( .A(n373), .B(n1621), .C(n370), .Z(n368) );
  CENX1 U1456 ( .A(n1564), .B(n236), .Z(product[26]) );
  CENX1 U1457 ( .A(n1657), .B(b[24]), .Z(n1366) );
  CIVX2 U1458 ( .A(n1585), .Z(n1657) );
  CNIVX1 U1459 ( .A(n1601), .Z(n1558) );
  CENX1 U1460 ( .A(n1667), .B(a[8]), .Z(n1601) );
  CIVX2 U1461 ( .A(n30), .Z(n1672) );
  CIVX2 U1462 ( .A(n1672), .Z(n1667) );
  CIVX2 U1463 ( .A(n87), .Z(n1700) );
  CIVDX1 U1464 ( .A(n55), .Z0(n1560), .Z1(n1561) );
  CIVX2 U1465 ( .A(n1575), .Z(n1676) );
  COR2X1 U1466 ( .A(n431), .B(n458), .Z(n1562) );
  COND2XL U1467 ( .A(n77), .B(n1201), .C(n1200), .D(n74), .Z(n922) );
  CENX1 U1468 ( .A(n1707), .B(n1703), .Z(n1158) );
  COND2X1 U1469 ( .A(n1158), .B(n100), .C(n102), .D(n1159), .Z(n884) );
  COND2XL U1470 ( .A(n91), .B(n1180), .C(n1179), .D(n89), .Z(n903) );
  CENX1 U1471 ( .A(n1664), .B(b[25]), .Z(n1334) );
  CENX1 U1472 ( .A(n1664), .B(n153), .Z(n1340) );
  CENX1 U1473 ( .A(n1658), .B(n156), .Z(n1368) );
  CENX1 U1474 ( .A(n1657), .B(n157), .Z(n1367) );
  CENX1 U1475 ( .A(n1684), .B(n1653), .Z(n1244) );
  CNIVXL U1476 ( .A(n120), .Z(n1708) );
  CNIVX2 U1477 ( .A(n120), .Z(n1707) );
  CEOX1 U1478 ( .A(a[12]), .B(n55), .Z(n1452) );
  CND2X1 U1479 ( .A(n1698), .B(a[22]), .Z(n1583) );
  COND2XL U1480 ( .A(n18), .B(n1362), .C(n1626), .D(n1361), .Z(n1076) );
  COND2XL U1481 ( .A(n18), .B(n1385), .C(n1626), .D(n1384), .Z(n1099) );
  COND2XL U1482 ( .A(n18), .B(n1363), .C(n1626), .D(n1362), .Z(n1077) );
  COND2XL U1483 ( .A(n18), .B(n1388), .C(n1626), .D(n1387), .Z(n1102) );
  CIVX1 U1484 ( .A(n292), .Z(n291) );
  COND2X1 U1485 ( .A(n77), .B(n1213), .C(n74), .D(n1212), .Z(n934) );
  CND2X2 U1486 ( .A(n1450), .B(n74), .Z(n77) );
  CENX1 U1487 ( .A(n1645), .B(n1690), .Z(n1212) );
  CND2X1 U1488 ( .A(n1600), .B(n394), .Z(n261) );
  CENX1 U1489 ( .A(n1668), .B(n1650), .Z(n1322) );
  CENXL U1490 ( .A(n1668), .B(n1651), .Z(n1321) );
  CIVX2 U1491 ( .A(n1683), .Z(n1681) );
  CEOX2 U1492 ( .A(a[18]), .B(n1693), .Z(n1449) );
  CENXL U1493 ( .A(n1692), .B(n1648), .Z(n1192) );
  CENXL U1494 ( .A(n1692), .B(n142), .Z(n1186) );
  CIVX1 U1495 ( .A(n71), .Z(n1691) );
  CENXL U1496 ( .A(n1687), .B(n1644), .Z(n1213) );
  CIVXL U1497 ( .A(n234), .Z(n389) );
  CIVX2 U1498 ( .A(n1560), .Z(n1684) );
  CANR1X1 U1499 ( .A(n390), .B(n241), .C(n238), .Z(n236) );
  CEOX4 U1500 ( .A(n1586), .B(a[4]), .Z(n1624) );
  CHA1XL U1501 ( .A(n853), .B(n892), .CO(n584), .S(n585) );
  COND2XL U1502 ( .A(n27), .B(n1341), .C(n24), .D(n1340), .Z(n1056) );
  CIVX1 U1503 ( .A(n229), .Z(n231) );
  CFA1XL U1504 ( .A(n943), .B(n1053), .CI(n1027), .CO(n554), .S(n555) );
  CFA1XL U1505 ( .A(n1003), .B(n584), .CI(n1111), .CO(n552), .S(n553) );
  COND2X1 U1506 ( .A(n91), .B(n1178), .C(n1177), .D(n89), .Z(n901) );
  CNR2XL U1507 ( .A(n85), .B(n1196), .Z(n1578) );
  CANR1X1 U1508 ( .A(n243), .B(n279), .C(n244), .Z(n1565) );
  CFA1XL U1509 ( .A(n955), .B(n993), .CI(n973), .CO(n776), .S(n777) );
  CANR1X1 U1510 ( .A(n221), .B(n241), .C(n222), .Z(n220) );
  CENXL U1511 ( .A(n1669), .B(n157), .Z(n1307) );
  CENXL U1512 ( .A(n1673), .B(n157), .Z(n1280) );
  CENXL U1513 ( .A(n1661), .B(n157), .Z(n1336) );
  CENXL U1514 ( .A(n1684), .B(n1648), .Z(n1249) );
  CENXL U1515 ( .A(n1684), .B(n1644), .Z(n1253) );
  CENXL U1516 ( .A(n1684), .B(n1651), .Z(n1246) );
  CENXL U1517 ( .A(n1684), .B(n146), .Z(n1241) );
  CENXL U1518 ( .A(n1684), .B(n142), .Z(n1243) );
  CENXL U1519 ( .A(n1684), .B(n1652), .Z(n1245) );
  CFA1XL U1520 ( .A(n1041), .B(n1095), .CI(n1067), .CO(n796), .S(n797) );
  CIVX1 U1521 ( .A(n330), .Z(n329) );
  CNIVX1 U1522 ( .A(n1006), .Z(n1563) );
  CENX1 U1523 ( .A(a[10]), .B(n1682), .Z(n1603) );
  COND2X1 U1524 ( .A(n69), .B(n1223), .C(n1222), .D(n66), .Z(n943) );
  CAN2X1 U1525 ( .A(n1562), .B(n1608), .Z(n1606) );
  CFA1XL U1526 ( .A(n915), .B(n1055), .CI(n945), .CO(n604), .S(n605) );
  CANR1X1 U1527 ( .A(n228), .B(n241), .C(n229), .Z(n227) );
  CND2X1 U1528 ( .A(n216), .B(n228), .Z(n214) );
  CNR2X1 U1529 ( .A(n234), .B(n239), .Z(n228) );
  CFA1XL U1530 ( .A(n952), .B(n1062), .CI(n1036), .CO(n732), .S(n733) );
  CNR2X1 U1531 ( .A(n295), .B(n298), .Z(n293) );
  CIVX1 U1532 ( .A(n295), .Z(n397) );
  COND2XL U1533 ( .A(n36), .B(n1306), .C(n1305), .D(n33), .Z(n1022) );
  COND2XL U1534 ( .A(n36), .B(n1308), .C(n1307), .D(n33), .Z(n1024) );
  COND2XL U1535 ( .A(n36), .B(n1328), .C(n1327), .D(n33), .Z(n1044) );
  COND2XL U1536 ( .A(n36), .B(n1307), .C(n1306), .D(n33), .Z(n1023) );
  COND2XL U1537 ( .A(n36), .B(n1310), .C(n1309), .D(n33), .Z(n1026) );
  COND2XL U1538 ( .A(n36), .B(n1330), .C(n33), .D(n1329), .Z(n1046) );
  COND2XL U1539 ( .A(n36), .B(n1671), .C(n1331), .D(n33), .Z(n862) );
  COND2XL U1540 ( .A(n36), .B(n1326), .C(n1325), .D(n33), .Z(n1042) );
  COND2XL U1541 ( .A(n36), .B(n1309), .C(n1308), .D(n33), .Z(n1025) );
  COND2XL U1542 ( .A(n36), .B(n1323), .C(n1322), .D(n33), .Z(n1039) );
  COND2XL U1543 ( .A(n36), .B(n1329), .C(n1328), .D(n33), .Z(n1045) );
  COND2XL U1544 ( .A(n36), .B(n1319), .C(n1318), .D(n33), .Z(n1035) );
  COND2XL U1545 ( .A(n36), .B(n1324), .C(n1323), .D(n33), .Z(n1040) );
  COND2XL U1546 ( .A(n36), .B(n1311), .C(n1310), .D(n33), .Z(n1027) );
  COND2XL U1547 ( .A(n36), .B(n1312), .C(n1311), .D(n33), .Z(n1028) );
  COND2XL U1548 ( .A(n36), .B(n1314), .C(n1313), .D(n33), .Z(n1030) );
  COND2XL U1549 ( .A(n36), .B(n1325), .C(n1324), .D(n33), .Z(n1041) );
  COND2XL U1550 ( .A(n36), .B(n1327), .C(n1326), .D(n33), .Z(n1043) );
  COND2X1 U1551 ( .A(n44), .B(n1285), .C(n1284), .D(n1559), .Z(n1002) );
  COND2XL U1552 ( .A(n69), .B(n1222), .C(n1221), .D(n66), .Z(n942) );
  CNR2IXL U1553 ( .B(n1706), .A(n66), .Z(n955) );
  COND2XL U1554 ( .A(n69), .B(n1221), .C(n1220), .D(n66), .Z(n941) );
  COND2XL U1555 ( .A(n69), .B(n1232), .C(n66), .D(n1231), .Z(n952) );
  COND2XL U1556 ( .A(n44), .B(n1281), .C(n1280), .D(n1559), .Z(n998) );
  COND2XL U1557 ( .A(n44), .B(n1282), .C(n1281), .D(n1559), .Z(n999) );
  COND2XL U1558 ( .A(n44), .B(n1283), .C(n1282), .D(n1559), .Z(n1000) );
  COND2XL U1559 ( .A(n44), .B(n1294), .C(n1293), .D(n1559), .Z(n1011) );
  COND2XL U1560 ( .A(n44), .B(n1680), .C(n1304), .D(n1559), .Z(n861) );
  COND2XL U1561 ( .A(n44), .B(n1301), .C(n1559), .D(n1300), .Z(n1018) );
  COND2XL U1562 ( .A(n44), .B(n1284), .C(n1283), .D(n1559), .Z(n1001) );
  COND2XL U1563 ( .A(n44), .B(n1289), .C(n1288), .D(n1559), .Z(n1006) );
  COND2XL U1564 ( .A(n44), .B(n1288), .C(n1287), .D(n1559), .Z(n1005) );
  COND2XL U1565 ( .A(n44), .B(n1298), .C(n1297), .D(n1559), .Z(n1015) );
  COND2XL U1566 ( .A(n44), .B(n1286), .C(n1285), .D(n1559), .Z(n1003) );
  COND2XL U1567 ( .A(n44), .B(n1303), .C(n1559), .D(n1302), .Z(n1020) );
  COND2XL U1568 ( .A(n44), .B(n1300), .C(n1299), .D(n1559), .Z(n1017) );
  COND2XL U1569 ( .A(n44), .B(n1292), .C(n1291), .D(n1559), .Z(n1009) );
  COND2XL U1570 ( .A(n44), .B(n1299), .C(n1298), .D(n1559), .Z(n1016) );
  COND2XL U1571 ( .A(n44), .B(n1295), .C(n1294), .D(n1559), .Z(n1012) );
  COND2XL U1572 ( .A(n44), .B(n1293), .C(n1292), .D(n1559), .Z(n1010) );
  CND2IX2 U1573 ( .B(n1602), .A(n1558), .Z(n44) );
  COND2X1 U1574 ( .A(n53), .B(n1270), .C(n1269), .D(n50), .Z(n988) );
  CFA1X1 U1575 ( .A(n936), .B(n1090), .CI(n990), .CO(n734), .S(n735) );
  COR2X1 U1576 ( .A(n671), .B(n688), .Z(n1611) );
  COND2X1 U1577 ( .A(n53), .B(n1265), .C(n1264), .D(n50), .Z(n983) );
  CND2X2 U1578 ( .A(n1583), .B(n1584), .Z(n95) );
  COND2XL U1579 ( .A(n1167), .B(n97), .C(n1166), .D(n95), .Z(n891) );
  COND2XL U1580 ( .A(n1167), .B(n95), .C(n1168), .D(n97), .Z(n892) );
  CENXL U1581 ( .A(n1657), .B(b[28]), .Z(n1362) );
  CENXL U1582 ( .A(n1684), .B(n153), .Z(n1236) );
  CIVX2 U1583 ( .A(n1585), .Z(n1659) );
  CENX2 U1584 ( .A(n1645), .B(n1694), .Z(n1195) );
  CIVX1 U1585 ( .A(n1697), .Z(n1694) );
  CIVX1 U1586 ( .A(n79), .Z(n1697) );
  COND1X1 U1587 ( .A(n330), .B(n313), .C(n314), .Z(n312) );
  CANR1X1 U1588 ( .A(n1614), .B(n321), .C(n316), .Z(n314) );
  CANR1X2 U1589 ( .A(n312), .B(n293), .C(n294), .Z(n292) );
  CIVX2 U1590 ( .A(n48), .Z(n1683) );
  COND1X2 U1591 ( .A(n245), .B(n262), .C(n246), .Z(n244) );
  CND2X4 U1592 ( .A(n89), .B(n1448), .Z(n91) );
  CENX4 U1593 ( .A(n1692), .B(a[20]), .Z(n89) );
  CENXL U1594 ( .A(n1686), .B(n148), .Z(n1219) );
  CENXL U1595 ( .A(n1676), .B(n148), .Z(n1288) );
  CENXL U1596 ( .A(n1684), .B(n148), .Z(n1240) );
  CENXL U1597 ( .A(n1664), .B(n148), .Z(n1344) );
  CENXL U1598 ( .A(n1657), .B(n148), .Z(n1375) );
  CENXL U1599 ( .A(n1669), .B(n148), .Z(n1315) );
  CHA1X1 U1600 ( .A(n854), .B(n904), .CO(n628), .S(n629) );
  COND2X1 U1601 ( .A(n97), .B(n1702), .C(n95), .D(n1171), .Z(n854) );
  CAN2XL U1602 ( .A(n389), .B(n235), .Z(n1564) );
  CNR2X1 U1603 ( .A(n218), .B(n223), .Z(n216) );
  CFA1XL U1604 ( .A(n901), .B(n961), .CI(n913), .CO(n558), .S(n559) );
  CENXL U1605 ( .A(n1640), .B(n1650), .Z(n1226) );
  CENXL U1606 ( .A(n1684), .B(n1650), .Z(n1247) );
  CENX4 U1607 ( .A(n1675), .B(a[10]), .Z(n50) );
  CIVX2 U1608 ( .A(n1679), .Z(n1675) );
  COND2X1 U1609 ( .A(n53), .B(n1263), .C(n1262), .D(n50), .Z(n981) );
  COND2X1 U1610 ( .A(n102), .B(n1704), .C(n100), .D(n1160), .Z(n853) );
  CENX4 U1611 ( .A(n1701), .B(a[24]), .Z(n100) );
  CENXL U1612 ( .A(n1667), .B(n1705), .Z(n1330) );
  CENXL U1613 ( .A(n1705), .B(n1695), .Z(n1198) );
  CENXL U1614 ( .A(n1705), .B(n1684), .Z(n1255) );
  COND1X1 U1615 ( .A(n352), .B(n340), .C(n341), .Z(n339) );
  CANR1X1 U1616 ( .A(n348), .B(n1618), .C(n343), .Z(n341) );
  CIVDX2 U1617 ( .A(n1660), .Z0(n1586), .Z1(n1585) );
  CIVX2 U1618 ( .A(n12), .Z(n1660) );
  CENXL U1619 ( .A(n1651), .B(n1701), .Z(n1161) );
  CENXL U1620 ( .A(n1644), .B(n1701), .Z(n1168) );
  COND1X2 U1621 ( .A(n280), .B(n292), .C(n281), .Z(n279) );
  CANR1X2 U1622 ( .A(n275), .B(n1600), .C(n268), .Z(n262) );
  CNIVX2 U1623 ( .A(n130), .Z(n1648) );
  COND1X1 U1624 ( .A(n299), .B(n295), .C(n296), .Z(n294) );
  CENXL U1625 ( .A(n1684), .B(n1649), .Z(n1248) );
  CENXL U1626 ( .A(n1674), .B(n1649), .Z(n1296) );
  CENX4 U1627 ( .A(n1685), .B(a[16]), .Z(n74) );
  CIVX4 U1628 ( .A(n1588), .Z(n1685) );
  CND2X1 U1629 ( .A(n1669), .B(n1654), .Z(n1567) );
  CND2X1 U1630 ( .A(n1671), .B(n1566), .Z(n1568) );
  CND2X1 U1631 ( .A(n1567), .B(n1568), .Z(n1317) );
  CIVXL U1632 ( .A(n1654), .Z(n1566) );
  CNIVX1 U1633 ( .A(n144), .Z(n1654) );
  COND2XL U1634 ( .A(n36), .B(n1318), .C(n1317), .D(n33), .Z(n1034) );
  CEOX1 U1635 ( .A(n619), .B(n638), .Z(n1569) );
  CEOX1 U1636 ( .A(n1569), .B(n636), .Z(n613) );
  CND2X1 U1637 ( .A(n636), .B(n638), .Z(n1570) );
  CND2X1 U1638 ( .A(n636), .B(n619), .Z(n1571) );
  CND2X1 U1639 ( .A(n638), .B(n619), .Z(n1572) );
  CND3X1 U1640 ( .A(n1570), .B(n1571), .C(n1572), .Z(n612) );
  CENXL U1641 ( .A(n1657), .B(n1646), .Z(n1386) );
  CENXL U1642 ( .A(n1662), .B(n1646), .Z(n1355) );
  CENXL U1643 ( .A(n1684), .B(n1646), .Z(n1251) );
  CENXL U1644 ( .A(n1640), .B(n1646), .Z(n1230) );
  CENXL U1645 ( .A(n1667), .B(n1646), .Z(n1326) );
  CENXL U1646 ( .A(n1687), .B(n1646), .Z(n1211) );
  CIVX8 U1647 ( .A(n1624), .Z(n24) );
  CENXL U1648 ( .A(n1587), .B(n151), .Z(n1217) );
  CENXL U1649 ( .A(n1684), .B(n151), .Z(n1238) );
  CENXL U1650 ( .A(n1678), .B(n151), .Z(n1286) );
  CENXL U1651 ( .A(n1670), .B(n151), .Z(n1313) );
  CENXL U1652 ( .A(n1659), .B(n151), .Z(n1373) );
  CENXL U1653 ( .A(n1664), .B(n151), .Z(n1342) );
  CENXL U1654 ( .A(n1681), .B(n151), .Z(n1261) );
  CANR1X2 U1655 ( .A(n257), .B(n1609), .C(n1610), .Z(n246) );
  COND2X1 U1656 ( .A(n1156), .B(n102), .C(n100), .D(n1155), .Z(n881) );
  CENXL U1657 ( .A(n1681), .B(n155), .Z(n1257) );
  CENXL U1658 ( .A(n1681), .B(n154), .Z(n1258) );
  CENXL U1659 ( .A(n1681), .B(n1651), .Z(n1269) );
  CIVXL U1660 ( .A(n1052), .Z(n1573) );
  CIVX1 U1661 ( .A(n1573), .Z(n1574) );
  CEOX2 U1662 ( .A(a[22]), .B(n1701), .Z(n1447) );
  CENXL U1663 ( .A(n1657), .B(b[26]), .Z(n1364) );
  CENXL U1664 ( .A(n1586), .B(b[29]), .Z(n1361) );
  CENXL U1665 ( .A(n1662), .B(n1645), .Z(n1356) );
  CENXL U1666 ( .A(n1645), .B(n1684), .Z(n1252) );
  CENXL U1667 ( .A(n1643), .B(n208), .Z(product[30]) );
  CANR1X1 U1668 ( .A(n1608), .B(n213), .C(n210), .Z(n208) );
  CENXL U1669 ( .A(n1642), .B(n199), .Z(product[31]) );
  CANR1X1 U1670 ( .A(n1606), .B(n1598), .C(n1605), .Z(n199) );
  CENXL U1671 ( .A(n1666), .B(b[25]), .Z(n1305) );
  CENXL U1672 ( .A(n1657), .B(b[25]), .Z(n1365) );
  CIVXL U1673 ( .A(n39), .Z(n1575) );
  CIVX2 U1674 ( .A(n39), .Z(n1679) );
  COR2XL U1675 ( .A(n53), .B(n1277), .Z(n1576) );
  COR2XL U1676 ( .A(n1276), .B(n50), .Z(n1577) );
  CND2X1 U1677 ( .A(n1576), .B(n1577), .Z(n995) );
  CENXL U1678 ( .A(n1681), .B(n1644), .Z(n1276) );
  CNR2XL U1679 ( .A(n82), .B(n1195), .Z(n1579) );
  CND2X2 U1680 ( .A(n1449), .B(n82), .Z(n85) );
  CENXL U1681 ( .A(n1692), .B(n1644), .Z(n1196) );
  CENX4 U1682 ( .A(n1687), .B(a[18]), .Z(n82) );
  CIVXL U1683 ( .A(n71), .Z(n1580) );
  CND2X1 U1684 ( .A(n1581), .B(n1582), .Z(n1584) );
  CIVX2 U1685 ( .A(n1698), .Z(n1581) );
  CIVXL U1686 ( .A(a[22]), .Z(n1582) );
  CNR2IXL U1687 ( .B(n1706), .A(n95), .Z(n895) );
  COND2XL U1688 ( .A(n97), .B(n1162), .C(n95), .D(n1161), .Z(n886) );
  CIVDX2 U1689 ( .A(n63), .Z0(n1588), .Z1(n1587) );
  CEO3X2 U1690 ( .A(n879), .B(n867), .C(n873), .Z(n457) );
  CND2XL U1691 ( .A(n879), .B(n873), .Z(n1589) );
  CND2XL U1692 ( .A(n879), .B(n867), .Z(n1590) );
  CND2XL U1693 ( .A(n873), .B(n867), .Z(n1591) );
  CND3XL U1694 ( .A(n1589), .B(n1590), .C(n1591), .Z(n456) );
  COR2X1 U1695 ( .A(n1154), .B(n102), .Z(n1592) );
  COR2XL U1696 ( .A(n1153), .B(n100), .Z(n1593) );
  CNR2IXL U1697 ( .B(n1706), .A(n114), .Z(n867) );
  COND2XL U1698 ( .A(n1147), .B(n107), .C(n105), .D(n1146), .Z(n873) );
  CENXL U1699 ( .A(n1647), .B(n1703), .Z(n1154) );
  CND2X4 U1700 ( .A(n100), .B(n1446), .Z(n102) );
  CND2XL U1701 ( .A(n433), .B(n460), .Z(n1595) );
  CND2X1 U1702 ( .A(n433), .B(n435), .Z(n1596) );
  CND2XL U1703 ( .A(n460), .B(n435), .Z(n1597) );
  CND2XL U1704 ( .A(n430), .B(n415), .Z(n198) );
  CENXL U1705 ( .A(n1648), .B(n1703), .Z(n1153) );
  CENXL U1706 ( .A(n1674), .B(n1648), .Z(n1297) );
  CENXL U1707 ( .A(n1687), .B(n1648), .Z(n1209) );
  CENXL U1708 ( .A(n1640), .B(n1648), .Z(n1228) );
  CENXL U1709 ( .A(n1684), .B(n1654), .Z(n1242) );
  COND2XL U1710 ( .A(n27), .B(n1337), .C(n24), .D(n1336), .Z(n1052) );
  CEOX2 U1711 ( .A(a[20]), .B(n1699), .Z(n1448) );
  COND1XL U1712 ( .A(n214), .B(n1565), .C(n215), .Z(n1598) );
  COND1XL U1713 ( .A(n214), .B(n242), .C(n215), .Z(n1599) );
  COND1XL U1714 ( .A(n214), .B(n1565), .C(n215), .Z(n213) );
  CNR2IXL U1715 ( .B(n1706), .A(n110), .Z(n871) );
  CIVX3 U1716 ( .A(a[0]), .Z(n6) );
  CIVXL U1717 ( .A(n312), .Z(n311) );
  CNIVX1 U1718 ( .A(n116), .Z(n1705) );
  CNIVX4 U1719 ( .A(n122), .Z(n1644) );
  CANR1X2 U1720 ( .A(n243), .B(n279), .C(n244), .Z(n242) );
  CNR2IXL U1721 ( .B(n1706), .A(n89), .Z(n907) );
  CENXL U1722 ( .A(n1688), .B(n148), .Z(n1200) );
  CEOXL U1723 ( .A(n186), .B(n338), .Z(product[11]) );
  CEOXL U1724 ( .A(n368), .B(n192), .Z(product[5]) );
  COND2X1 U1725 ( .A(n18), .B(n1387), .C(n1626), .D(n1386), .Z(n1101) );
  CNR2IXL U1726 ( .B(n1706), .A(n33), .Z(n1047) );
  COND2X1 U1727 ( .A(n18), .B(n1382), .C(n1626), .D(n1381), .Z(n1096) );
  CENX1 U1728 ( .A(n1685), .B(n1653), .Z(n1223) );
  CENX1 U1729 ( .A(n1685), .B(n1652), .Z(n1224) );
  COND2X1 U1730 ( .A(n77), .B(n1212), .C(n1211), .D(n74), .Z(n933) );
  CNR2IXL U1731 ( .B(n1706), .A(n1559), .Z(n1021) );
  CEOXL U1732 ( .A(n376), .B(n194), .Z(product[3]) );
  CNIVX1 U1733 ( .A(n134), .Z(n1650) );
  CNIVX2 U1734 ( .A(n138), .Z(n1652) );
  CNIVX1 U1735 ( .A(n140), .Z(n1653) );
  CANR1X1 U1736 ( .A(n229), .B(n216), .C(n217), .Z(n215) );
  CEOXL U1737 ( .A(n170), .B(n227), .Z(product[27]) );
  CND2XL U1738 ( .A(n388), .B(n226), .Z(n170) );
  CEOXL U1739 ( .A(n220), .B(n169), .Z(product[28]) );
  CND2XL U1740 ( .A(n387), .B(n219), .Z(n169) );
  CND2XL U1741 ( .A(n263), .B(n1607), .Z(n252) );
  CND2XL U1742 ( .A(n320), .B(n1614), .Z(n313) );
  CND2XL U1743 ( .A(n397), .B(n296), .Z(n179) );
  CIVX1 U1744 ( .A(n303), .Z(n301) );
  CEOXL U1745 ( .A(n182), .B(n319), .Z(product[15]) );
  CND2XL U1746 ( .A(n1614), .B(n318), .Z(n182) );
  CEOXL U1747 ( .A(n177), .B(n286), .Z(product[20]) );
  CND2XL U1748 ( .A(n1611), .B(n285), .Z(n177) );
  CEOXL U1749 ( .A(n176), .B(n278), .Z(product[21]) );
  CND2XL U1750 ( .A(n394), .B(n273), .Z(n176) );
  CEOXL U1751 ( .A(n181), .B(n311), .Z(product[16]) );
  CND2XL U1752 ( .A(n399), .B(n306), .Z(n181) );
  CND2XL U1753 ( .A(n1612), .B(n303), .Z(n180) );
  CND2XL U1754 ( .A(n1613), .B(n290), .Z(n178) );
  CND2XL U1755 ( .A(n1612), .B(n399), .Z(n298) );
  CIVX1 U1756 ( .A(n270), .Z(n268) );
  CANR1X1 U1757 ( .A(n1616), .B(n357), .C(n354), .Z(n352) );
  CNR2XL U1758 ( .A(n322), .B(n327), .Z(n320) );
  CND2XL U1759 ( .A(n1618), .B(n345), .Z(n187) );
  CND2XL U1760 ( .A(n404), .B(n337), .Z(n186) );
  CND2XL U1761 ( .A(n1616), .B(n356), .Z(n189) );
  CND2XL U1762 ( .A(n1617), .B(n350), .Z(n188) );
  CND2XL U1763 ( .A(n402), .B(n328), .Z(n184) );
  COR2X1 U1764 ( .A(n1631), .B(n650), .Z(n1600) );
  CND2XL U1765 ( .A(n767), .B(n778), .Z(n323) );
  COND1X1 U1766 ( .A(n358), .B(n360), .C(n359), .Z(n357) );
  CANR1X1 U1767 ( .A(n365), .B(n1620), .C(n362), .Z(n360) );
  CND2XL U1768 ( .A(n791), .B(n800), .Z(n334) );
  COR2XL U1769 ( .A(n819), .B(n826), .Z(n1617) );
  CND2XL U1770 ( .A(n1620), .B(n364), .Z(n191) );
  CND2XL U1771 ( .A(n410), .B(n367), .Z(n192) );
  CND2XL U1772 ( .A(n849), .B(n864), .Z(n375) );
  CND2XL U1773 ( .A(n833), .B(n838), .Z(n359) );
  CEO3X1 U1774 ( .A(n434), .B(n416), .C(n432), .Z(n415) );
  CEO3X1 U1775 ( .A(n436), .B(n418), .C(n417), .Z(n416) );
  CEO3X1 U1776 ( .A(n420), .B(n438), .C(n419), .Z(n417) );
  COR2XL U1777 ( .A(n1135), .B(n1105), .Z(n1622) );
  COND2X1 U1778 ( .A(n1158), .B(n102), .C(n100), .D(n1157), .Z(n883) );
  CND2IXL U1779 ( .B(n1706), .A(n1681), .Z(n1279) );
  CND2XL U1780 ( .A(n412), .B(n375), .Z(n194) );
  CENX4 U1781 ( .A(n1561), .B(a[14]), .Z(n66) );
  CND2X4 U1782 ( .A(n1457), .B(n1626), .Z(n18) );
  CEOX2 U1783 ( .A(a[2]), .B(n1659), .Z(n1457) );
  CENX1 U1784 ( .A(a[8]), .B(n1676), .Z(n1602) );
  CNIVX1 U1785 ( .A(n132), .Z(n1649) );
  CNIVX1 U1786 ( .A(n136), .Z(n1651) );
  CND2IX2 U1787 ( .B(n1603), .A(n50), .Z(n53) );
  CND2X4 U1788 ( .A(n1451), .B(n66), .Z(n69) );
  CEOX2 U1789 ( .A(a[14]), .B(n1587), .Z(n1451) );
  CNIVX1 U1790 ( .A(n126), .Z(n1646) );
  CEOXL U1791 ( .A(a[28]), .B(n109), .Z(n1444) );
  CEOXL U1792 ( .A(a[30]), .B(n113), .Z(n1443) );
  CND2XL U1793 ( .A(n1622), .B(n380), .Z(n195) );
  CENX1 U1794 ( .A(n260), .B(n174), .Z(product[23]) );
  CND2X1 U1795 ( .A(n1607), .B(n259), .Z(n174) );
  CENX1 U1796 ( .A(n241), .B(n172), .Z(product[25]) );
  CEOXL U1797 ( .A(n1599), .B(n1604), .Z(product[29]) );
  CAN2XL U1798 ( .A(n1608), .B(n212), .Z(n1604) );
  COND1XL U1799 ( .A(n223), .B(n231), .C(n226), .Z(n222) );
  CANR1XL U1800 ( .A(n1607), .B(n264), .C(n257), .Z(n253) );
  COND1XL U1801 ( .A(n252), .B(n278), .C(n253), .Z(n251) );
  CNR2IXL U1802 ( .B(n228), .A(n223), .Z(n221) );
  CAOR1X1 U1803 ( .A(n210), .B(n1562), .C(n205), .Z(n1605) );
  CND2X1 U1804 ( .A(n1611), .B(n1613), .Z(n280) );
  CNR2X1 U1805 ( .A(n563), .B(n586), .Z(n239) );
  CENX1 U1806 ( .A(n297), .B(n179), .Z(product[18]) );
  CENX1 U1807 ( .A(n271), .B(n175), .Z(product[22]) );
  CND2X1 U1808 ( .A(n1600), .B(n270), .Z(n175) );
  COND1XL U1809 ( .A(n272), .B(n278), .C(n273), .Z(n271) );
  CENX1 U1810 ( .A(n304), .B(n180), .Z(product[17]) );
  COND1XL U1811 ( .A(n305), .B(n311), .C(n306), .Z(n304) );
  CENX1 U1812 ( .A(n291), .B(n178), .Z(product[19]) );
  CNR2X2 U1813 ( .A(n539), .B(n562), .Z(n234) );
  COR2X1 U1814 ( .A(n609), .B(n630), .Z(n1607) );
  CANR1XL U1815 ( .A(n1613), .B(n291), .C(n288), .Z(n286) );
  CEOX1 U1816 ( .A(n183), .B(n324), .Z(product[14]) );
  CND2X1 U1817 ( .A(n401), .B(n323), .Z(n183) );
  CANR1XL U1818 ( .A(n402), .B(n329), .C(n326), .Z(n324) );
  CANR1XL U1819 ( .A(n320), .B(n329), .C(n321), .Z(n319) );
  COR2X1 U1820 ( .A(n459), .B(n486), .Z(n1608) );
  CND2X1 U1821 ( .A(n539), .B(n562), .Z(n235) );
  CND2X1 U1822 ( .A(n513), .B(n538), .Z(n226) );
  CND2X1 U1823 ( .A(n609), .B(n630), .Z(n259) );
  CND2X1 U1824 ( .A(n487), .B(n512), .Z(n219) );
  COR2X1 U1825 ( .A(n587), .B(n608), .Z(n1609) );
  CAN2X1 U1826 ( .A(n587), .B(n608), .Z(n1610) );
  CND2X1 U1827 ( .A(n1618), .B(n1617), .Z(n340) );
  CANR1X1 U1828 ( .A(n331), .B(n339), .C(n332), .Z(n330) );
  CNR2X1 U1829 ( .A(n333), .B(n336), .Z(n331) );
  COND1XL U1830 ( .A(n337), .B(n333), .C(n334), .Z(n332) );
  CENX1 U1831 ( .A(n189), .B(n357), .Z(product[8]) );
  COND1XL U1832 ( .A(n328), .B(n322), .C(n323), .Z(n321) );
  CENX1 U1833 ( .A(n335), .B(n185), .Z(product[12]) );
  CND2X1 U1834 ( .A(n403), .B(n334), .Z(n185) );
  COND1XL U1835 ( .A(n336), .B(n338), .C(n337), .Z(n335) );
  CENX1 U1836 ( .A(n188), .B(n351), .Z(product[9]) );
  CENX1 U1837 ( .A(n329), .B(n184), .Z(product[13]) );
  CNR2X1 U1838 ( .A(n767), .B(n778), .Z(n322) );
  CNR2X1 U1839 ( .A(n739), .B(n752), .Z(n305) );
  CEOX1 U1840 ( .A(n346), .B(n187), .Z(product[10]) );
  CANR1XL U1841 ( .A(n1617), .B(n351), .C(n348), .Z(n346) );
  COR2X1 U1842 ( .A(n723), .B(n738), .Z(n1612) );
  COR2X1 U1843 ( .A(n689), .B(n706), .Z(n1613) );
  CND2X1 U1844 ( .A(n651), .B(n670), .Z(n273) );
  CND2X1 U1845 ( .A(n739), .B(n752), .Z(n306) );
  CND2X1 U1846 ( .A(n707), .B(n722), .Z(n296) );
  COR2X1 U1847 ( .A(n753), .B(n766), .Z(n1614) );
  CND2X1 U1848 ( .A(n689), .B(n706), .Z(n290) );
  CND2X1 U1849 ( .A(n631), .B(n650), .Z(n270) );
  CND2X1 U1850 ( .A(n671), .B(n688), .Z(n285) );
  CND2X1 U1851 ( .A(n723), .B(n738), .Z(n303) );
  CND2X1 U1852 ( .A(n753), .B(n766), .Z(n318) );
  COND1XL U1853 ( .A(n368), .B(n366), .C(n367), .Z(n365) );
  CAN2X1 U1854 ( .A(n1619), .B(n198), .Z(n1642) );
  CND3XL U1855 ( .A(n1634), .B(n1635), .C(n1636), .Z(n650) );
  CNR2X1 U1856 ( .A(n801), .B(n810), .Z(n336) );
  CNR2X1 U1857 ( .A(n791), .B(n800), .Z(n333) );
  CENX1 U1858 ( .A(n1615), .B(n653), .Z(n651) );
  CENX1 U1859 ( .A(n655), .B(n672), .Z(n1615) );
  CNR2X1 U1860 ( .A(n779), .B(n790), .Z(n327) );
  COR2X1 U1861 ( .A(n827), .B(n832), .Z(n1616) );
  CND2X1 U1862 ( .A(n779), .B(n790), .Z(n328) );
  COR2X1 U1863 ( .A(n811), .B(n818), .Z(n1618) );
  CND2X1 U1864 ( .A(n801), .B(n810), .Z(n337) );
  CND2X1 U1865 ( .A(n819), .B(n826), .Z(n350) );
  CND2X1 U1866 ( .A(n827), .B(n832), .Z(n356) );
  CND2X1 U1867 ( .A(n811), .B(n818), .Z(n345) );
  COR2X1 U1868 ( .A(n430), .B(n415), .Z(n1619) );
  CENX1 U1869 ( .A(n191), .B(n365), .Z(product[6]) );
  CEOXL U1870 ( .A(n360), .B(n190), .Z(product[7]) );
  CND2X1 U1871 ( .A(n408), .B(n359), .Z(n190) );
  CNR2X1 U1872 ( .A(n833), .B(n838), .Z(n358) );
  CNR2X1 U1873 ( .A(n843), .B(n846), .Z(n366) );
  CNR2X1 U1874 ( .A(n849), .B(n864), .Z(n374) );
  COR2X1 U1875 ( .A(n839), .B(n842), .Z(n1620) );
  CND2X1 U1876 ( .A(n843), .B(n846), .Z(n367) );
  CND2X1 U1877 ( .A(n839), .B(n842), .Z(n364) );
  CND2X1 U1878 ( .A(n847), .B(n848), .Z(n372) );
  CND2X1 U1879 ( .A(n1135), .B(n1105), .Z(n380) );
  COR2X1 U1880 ( .A(n847), .B(n848), .Z(n1621) );
  CENX1 U1881 ( .A(n193), .B(n373), .Z(product[4]) );
  CND2XL U1882 ( .A(n1621), .B(n372), .Z(n193) );
  CENX1 U1883 ( .A(n1653), .B(n1689), .Z(n1204) );
  CENX1 U1884 ( .A(n1688), .B(n1652), .Z(n1205) );
  CENX1 U1885 ( .A(n1666), .B(n155), .Z(n1309) );
  CENX1 U1886 ( .A(n1673), .B(n155), .Z(n1282) );
  CENX1 U1887 ( .A(n1657), .B(n155), .Z(n1369) );
  CENX1 U1888 ( .A(n1707), .B(n1684), .Z(n1254) );
  CENX1 U1889 ( .A(n1663), .B(n1652), .Z(n1349) );
  CENX1 U1890 ( .A(n1664), .B(n1653), .Z(n1348) );
  CENX1 U1891 ( .A(n1707), .B(n1587), .Z(n1233) );
  CENX1 U1892 ( .A(n1707), .B(n1699), .Z(n1182) );
  CENX1 U1893 ( .A(n1657), .B(n1644), .Z(n1388) );
  CENX1 U1894 ( .A(n1707), .B(n1662), .Z(n1358) );
  CENX1 U1895 ( .A(n1657), .B(n1648), .Z(n1384) );
  CENX1 U1896 ( .A(n1707), .B(n1670), .Z(n1329) );
  CENX1 U1897 ( .A(n1663), .B(n1651), .Z(n1350) );
  CENX1 U1898 ( .A(n1653), .B(n1699), .Z(n1172) );
  CENX1 U1899 ( .A(n1647), .B(n1686), .Z(n1229) );
  CENX1 U1900 ( .A(n1707), .B(n1695), .Z(n1197) );
  CIVX2 U1901 ( .A(n1700), .Z(n1698) );
  CIVX2 U1902 ( .A(n1683), .Z(n1682) );
  CIVX2 U1903 ( .A(n1700), .Z(n1699) );
  CENX1 U1904 ( .A(n1651), .B(n1695), .Z(n1189) );
  CENX1 U1905 ( .A(n1653), .B(n1695), .Z(n1187) );
  CENX1 U1906 ( .A(n1647), .B(n1694), .Z(n1193) );
  CENX1 U1907 ( .A(n1586), .B(n1651), .Z(n1381) );
  CNR2IX1 U1908 ( .B(n1706), .A(n1626), .Z(n1105) );
  CENX1 U1909 ( .A(n1698), .B(n1648), .Z(n1177) );
  CENX1 U1910 ( .A(n1699), .B(n1644), .Z(n1181) );
  CENX1 U1911 ( .A(n1676), .B(n1653), .Z(n1292) );
  CENX1 U1912 ( .A(n1669), .B(n1653), .Z(n1319) );
  CENX1 U1913 ( .A(n1676), .B(n1652), .Z(n1293) );
  CENX1 U1914 ( .A(n1667), .B(n1647), .Z(n1325) );
  CENX1 U1915 ( .A(n1647), .B(n1678), .Z(n1298) );
  CENX1 U1916 ( .A(n1666), .B(n1652), .Z(n1320) );
  CENX1 U1917 ( .A(n1698), .B(n1652), .Z(n1173) );
  CENX1 U1918 ( .A(n1667), .B(n1644), .Z(n1328) );
  CENX1 U1919 ( .A(n1675), .B(n1651), .Z(n1294) );
  CENX1 U1920 ( .A(n1666), .B(n1648), .Z(n1324) );
  CENX1 U1921 ( .A(n1662), .B(n1644), .Z(n1357) );
  CENX1 U1922 ( .A(n1647), .B(n1684), .Z(n1250) );
  CENX1 U1923 ( .A(n1658), .B(n1647), .Z(n1385) );
  CENX1 U1924 ( .A(n1651), .B(n1699), .Z(n1174) );
  CENX1 U1925 ( .A(n1658), .B(n1652), .Z(n1380) );
  CENX1 U1926 ( .A(n1658), .B(n1653), .Z(n1379) );
  CENX1 U1927 ( .A(n1662), .B(n1647), .Z(n1354) );
  CENX1 U1928 ( .A(n1664), .B(n1648), .Z(n1353) );
  CENX1 U1929 ( .A(n1685), .B(n1651), .Z(n1225) );
  CENX1 U1930 ( .A(n1693), .B(n1652), .Z(n1188) );
  CENX1 U1931 ( .A(n1644), .B(n1703), .Z(n1157) );
  CENX1 U1932 ( .A(n1662), .B(n1706), .Z(n1359) );
  CNR2IX1 U1933 ( .B(n1706), .A(n24), .Z(n1075) );
  CENX1 U1934 ( .A(n1586), .B(n1706), .Z(n1390) );
  CNR2IXL U1935 ( .B(n1706), .A(n58), .Z(n975) );
  CNR2IX1 U1936 ( .B(n1706), .A(n74), .Z(n937) );
  CNR2IXL U1937 ( .B(n1706), .A(n105), .Z(n877) );
  CND2X1 U1938 ( .A(n1449), .B(n82), .Z(n1633) );
  CNIVX1 U1939 ( .A(n980), .Z(n1629) );
  CEOX1 U1940 ( .A(n850), .B(n878), .Z(n429) );
  CNR2IX1 U1941 ( .B(n1706), .A(n6), .Z(product[0]) );
  CENX1 U1942 ( .A(n1677), .B(n146), .Z(n1289) );
  CENX1 U1943 ( .A(n1668), .B(n146), .Z(n1316) );
  CENX1 U1944 ( .A(n1688), .B(n142), .Z(n1203) );
  CENX1 U1945 ( .A(n1689), .B(n146), .Z(n1201) );
  CENX1 U1946 ( .A(n1673), .B(n156), .Z(n1281) );
  CENX1 U1947 ( .A(n1661), .B(n156), .Z(n1337) );
  CENX1 U1948 ( .A(n1658), .B(n152), .Z(n1372) );
  CENX1 U1949 ( .A(n1664), .B(n142), .Z(n1347) );
  CENX1 U1950 ( .A(n1657), .B(n146), .Z(n1376) );
  CENX1 U1951 ( .A(n1657), .B(n154), .Z(n1370) );
  CENX1 U1952 ( .A(n1708), .B(n109), .Z(n1142) );
  CENX1 U1953 ( .A(n104), .B(a[28]), .Z(n110) );
  CENX1 U1954 ( .A(n1662), .B(b[27]), .Z(n1332) );
  CENX1 U1955 ( .A(n1708), .B(n113), .Z(n1137) );
  CENX1 U1956 ( .A(n109), .B(a[30]), .Z(n114) );
  CENX1 U1957 ( .A(n1661), .B(n154), .Z(n1339) );
  CENX1 U1958 ( .A(n1658), .B(n142), .Z(n1378) );
  CENX1 U1959 ( .A(n1587), .B(n150), .Z(n1218) );
  CENX1 U1960 ( .A(n1647), .B(n104), .Z(n1145) );
  CENX1 U1961 ( .A(n1686), .B(n142), .Z(n1222) );
  CENX1 U1962 ( .A(n1669), .B(n150), .Z(n1314) );
  CENX1 U1963 ( .A(n1676), .B(n142), .Z(n1291) );
  CENX1 U1964 ( .A(n1666), .B(n142), .Z(n1318) );
  CENX1 U1965 ( .A(n1666), .B(n154), .Z(n1310) );
  CENX1 U1966 ( .A(n1675), .B(n154), .Z(n1283) );
  CENX1 U1967 ( .A(n1669), .B(n156), .Z(n1308) );
  CENX1 U1968 ( .A(n1684), .B(n150), .Z(n1239) );
  CENX1 U1969 ( .A(n1669), .B(b[24]), .Z(n1306) );
  CENXL U1970 ( .A(n1644), .B(n104), .Z(n1148) );
  CENX1 U1971 ( .A(n1644), .B(n109), .Z(n1141) );
  CENX1 U1972 ( .A(n1664), .B(n146), .Z(n1345) );
  CENX1 U1973 ( .A(n1664), .B(n150), .Z(n1343) );
  CENX1 U1974 ( .A(n1686), .B(n146), .Z(n1220) );
  CND2X1 U1975 ( .A(n1444), .B(n110), .Z(n112) );
  CND2X1 U1976 ( .A(n1443), .B(n114), .Z(n115) );
  CNIVXL U1980 ( .A(n63), .Z(n1640) );
  COND2XL U1981 ( .A(n18), .B(n1585), .C(n1391), .D(n1626), .Z(n864) );
  CIVX1 U1982 ( .A(n1054), .Z(n1627) );
  CIVX2 U1983 ( .A(n1627), .Z(n1628) );
  CIVX1 U1984 ( .A(n1672), .Z(n1670) );
  CIVX1 U1985 ( .A(n1672), .Z(n1669) );
  CEO3XL U1986 ( .A(n635), .B(n652), .C(n633), .Z(n1631) );
  CIVX2 U1987 ( .A(n242), .Z(n241) );
  CENX1 U1988 ( .A(n1708), .B(n104), .Z(n1149) );
  CIVXL U1989 ( .A(n218), .Z(n387) );
  COND1X1 U1990 ( .A(n226), .B(n218), .C(n219), .Z(n217) );
  CNR2X2 U1991 ( .A(n487), .B(n512), .Z(n218) );
  CENX1 U1992 ( .A(n1640), .B(n1644), .Z(n1232) );
  CND2IXL U1993 ( .B(n1706), .A(n1640), .Z(n1235) );
  CIVX2 U1994 ( .A(n1580), .Z(n1689) );
  CIVX2 U1995 ( .A(n1691), .Z(n1687) );
  COND2XL U1996 ( .A(n69), .B(n1218), .C(n1217), .D(n66), .Z(n938) );
  COND2XL U1997 ( .A(n69), .B(n1219), .C(n1218), .D(n66), .Z(n939) );
  COND2XL U1998 ( .A(n69), .B(n1220), .C(n1219), .D(n66), .Z(n940) );
  COND2XL U1999 ( .A(n69), .B(n1230), .C(n66), .D(n1229), .Z(n950) );
  COND2XL U2000 ( .A(n69), .B(n1226), .C(n1225), .D(n66), .Z(n946) );
  CIVX2 U2001 ( .A(n1696), .Z(n1692) );
  CENX1 U2002 ( .A(n1657), .B(n1654), .Z(n1377) );
  CENX1 U2003 ( .A(n251), .B(n173), .Z(product[24]) );
  CIVXL U2004 ( .A(n1610), .Z(n1632) );
  CIVX1 U2005 ( .A(n1585), .Z(n1658) );
  COND2XL U2006 ( .A(n18), .B(n1378), .C(n1626), .D(n1377), .Z(n1092) );
  COND2XL U2007 ( .A(n1152), .B(n100), .C(n1153), .D(n102), .Z(n878) );
  COND2XL U2008 ( .A(n1154), .B(n100), .C(n1155), .D(n102), .Z(n880) );
  COND2XL U2009 ( .A(n1156), .B(n100), .C(n1157), .D(n102), .Z(n882) );
  CNR2IXL U2010 ( .B(n1706), .A(n100), .Z(n885) );
  CND2IXL U2011 ( .B(n1706), .A(n1701), .Z(n1171) );
  CIVXL U2012 ( .A(n1691), .Z(n1690) );
  CENX1 U2013 ( .A(n1654), .B(n1689), .Z(n1202) );
  CENX1 U2014 ( .A(n1651), .B(n1690), .Z(n1206) );
  CENX1 U2015 ( .A(n1647), .B(n1690), .Z(n1210) );
  CND2XL U2016 ( .A(n653), .B(n672), .Z(n1634) );
  CND2XL U2017 ( .A(n653), .B(n655), .Z(n1635) );
  CND2X1 U2018 ( .A(n672), .B(n655), .Z(n1636) );
  CEO3X1 U2019 ( .A(n920), .B(n934), .C(n1060), .Z(n703) );
  CND2XL U2020 ( .A(n920), .B(n1060), .Z(n1637) );
  CND2XL U2021 ( .A(n920), .B(n934), .Z(n1638) );
  CND2XL U2022 ( .A(n1060), .B(n934), .Z(n1639) );
  COND2XL U2023 ( .A(n53), .B(n1258), .C(n1257), .D(n50), .Z(n976) );
  COND2XL U2024 ( .A(n53), .B(n1259), .C(n1258), .D(n50), .Z(n977) );
  COND2XL U2025 ( .A(n53), .B(n1274), .C(n50), .D(n1273), .Z(n992) );
  COND2XL U2026 ( .A(n53), .B(n1260), .C(n1259), .D(n50), .Z(n978) );
  CNR2IXL U2027 ( .B(n1706), .A(n50), .Z(n997) );
  COND2XL U2028 ( .A(n53), .B(n1261), .C(n1260), .D(n50), .Z(n979) );
  COND2XL U2029 ( .A(n53), .B(n1268), .C(n1267), .D(n50), .Z(n986) );
  COND2XL U2030 ( .A(n53), .B(n1271), .C(n1270), .D(n50), .Z(n989) );
  COND2XL U2031 ( .A(n53), .B(n1266), .C(n1265), .D(n50), .Z(n984) );
  COND2XL U2032 ( .A(n53), .B(n1269), .C(n1268), .D(n50), .Z(n987) );
  COND2XL U2033 ( .A(n53), .B(n1278), .C(n50), .D(n1277), .Z(n996) );
  COND2XL U2034 ( .A(n53), .B(n1272), .C(n1271), .D(n50), .Z(n990) );
  COND2XL U2035 ( .A(n53), .B(n1683), .C(n1279), .D(n50), .Z(n860) );
  COND2XL U2036 ( .A(n53), .B(n1276), .C(n50), .D(n1275), .Z(n994) );
  COND2XL U2037 ( .A(n53), .B(n1275), .C(n1274), .D(n50), .Z(n993) );
  COND2XL U2038 ( .A(n53), .B(n1262), .C(n1261), .D(n50), .Z(n980) );
  CNR2X1 U2039 ( .A(n651), .B(n670), .Z(n272) );
  CENX1 U2040 ( .A(n1647), .B(n1699), .Z(n1178) );
  COND2XL U2041 ( .A(n27), .B(n1339), .C(n24), .D(n1338), .Z(n1054) );
  CENXL U2042 ( .A(n1661), .B(n155), .Z(n1338) );
  COND2X1 U2043 ( .A(n1633), .B(n1197), .C(n82), .D(n1196), .Z(n919) );
  COND1X2 U2044 ( .A(n240), .B(n234), .C(n235), .Z(n229) );
  CND2IXL U2045 ( .B(n1706), .A(n1657), .Z(n1391) );
  CENXL U2046 ( .A(n1677), .B(n152), .Z(n1285) );
  CNR2X1 U2047 ( .A(n245), .B(n261), .Z(n243) );
  COND2XL U2048 ( .A(n69), .B(n1588), .C(n1235), .D(n66), .Z(n858) );
  CIVX1 U2049 ( .A(n1588), .Z(n1686) );
  CENX1 U2050 ( .A(n1654), .B(n1694), .Z(n1185) );
  CND2IXL U2051 ( .B(n1706), .A(n1661), .Z(n1360) );
  CND2IXL U2052 ( .B(n1706), .A(n1673), .Z(n1304) );
  CENX1 U2053 ( .A(n1674), .B(n1644), .Z(n1301) );
  COND1XL U2054 ( .A(n261), .B(n278), .C(n262), .Z(n260) );
  COND1XL U2055 ( .A(n298), .B(n311), .C(n299), .Z(n297) );
  COND2XL U2056 ( .A(n77), .B(n1691), .C(n1216), .D(n74), .Z(n857) );
  CEOX1 U2057 ( .A(a[16]), .B(n1689), .Z(n1450) );
  CIVX2 U2058 ( .A(n1697), .Z(n1693) );
  CIVXL U2059 ( .A(n262), .Z(n264) );
  CNIVX4 U2060 ( .A(n124), .Z(n1645) );
  CIVX1 U2061 ( .A(n1671), .Z(n1666) );
  CIVXL U2062 ( .A(n1694), .Z(n1641) );
  CND2X1 U2063 ( .A(n563), .B(n586), .Z(n240) );
  CND2XL U2064 ( .A(n390), .B(n240), .Z(n172) );
  CIVX1 U2065 ( .A(n240), .Z(n238) );
  CND2XL U2066 ( .A(n1609), .B(n1632), .Z(n173) );
  CAN2XL U2067 ( .A(n1562), .B(n207), .Z(n1643) );
  CND2X1 U2068 ( .A(n1609), .B(n1607), .Z(n245) );
  COND2XL U2069 ( .A(n1633), .B(n1186), .C(n82), .D(n1185), .Z(n908) );
  COND2XL U2070 ( .A(n1633), .B(n1189), .C(n1188), .D(n82), .Z(n911) );
  CNR2IXL U2071 ( .B(n1706), .A(n82), .Z(n921) );
  COND2XL U2072 ( .A(n1633), .B(n1188), .C(n82), .D(n1187), .Z(n910) );
  COND2XL U2073 ( .A(n1633), .B(n1187), .C(n1186), .D(n82), .Z(n909) );
  COND2XL U2074 ( .A(n1633), .B(n1194), .C(n82), .D(n1193), .Z(n916) );
  COND2XL U2075 ( .A(n1633), .B(n1641), .C(n1199), .D(n82), .Z(n856) );
  COND2XL U2076 ( .A(n85), .B(n1191), .C(n1190), .D(n82), .Z(n913) );
  COND2XL U2077 ( .A(n85), .B(n1190), .C(n82), .D(n1189), .Z(n912) );
  COND2XL U2078 ( .A(n1633), .B(n1198), .C(n82), .D(n1197), .Z(n920) );
  COND2XL U2079 ( .A(n1633), .B(n1193), .C(n1192), .D(n82), .Z(n915) );
  COND2XL U2080 ( .A(n85), .B(n1195), .C(n1194), .D(n82), .Z(n917) );
  CND2IXL U2081 ( .B(n1706), .A(n1687), .Z(n1216) );
  CIVX4 U2082 ( .A(n1702), .Z(n1701) );
  CND2X4 U2083 ( .A(n1456), .B(n24), .Z(n27) );
  CENX4 U2084 ( .A(n1682), .B(a[12]), .Z(n58) );
  CND2X4 U2085 ( .A(n1452), .B(n58), .Z(n61) );
  CIVXL U2086 ( .A(n1665), .Z(n1661) );
  CIVXL U2087 ( .A(n1672), .Z(n1668) );
  CIVXL U2088 ( .A(n30), .Z(n1671) );
  CIVXL U2089 ( .A(n1680), .Z(n1673) );
  CIVXL U2090 ( .A(n1680), .Z(n1674) );
  CIVXL U2091 ( .A(n1575), .Z(n1677) );
  CIVXL U2092 ( .A(n1680), .Z(n1678) );
  CIVXL U2093 ( .A(n39), .Z(n1680) );
  CIVXL U2094 ( .A(n1691), .Z(n1688) );
  CIVXL U2095 ( .A(n1697), .Z(n1695) );
  CIVXL U2096 ( .A(n79), .Z(n1696) );
  CIVX1 U2097 ( .A(n93), .Z(n1702) );
  CIVX1 U2098 ( .A(n99), .Z(n1704) );
  CIVX2 U2099 ( .A(n374), .Z(n412) );
  CIVX2 U2100 ( .A(n366), .Z(n410) );
  CIVX2 U2101 ( .A(n358), .Z(n408) );
  CIVX2 U2102 ( .A(n336), .Z(n404) );
  CIVX2 U2103 ( .A(n333), .Z(n403) );
  CIVX2 U2104 ( .A(n322), .Z(n401) );
  CIVX2 U2105 ( .A(n223), .Z(n388) );
  CIVX2 U2106 ( .A(n380), .Z(n378) );
  CIVX2 U2107 ( .A(n372), .Z(n370) );
  CIVX2 U2108 ( .A(n364), .Z(n362) );
  CIVX2 U2109 ( .A(n356), .Z(n354) );
  CIVX2 U2110 ( .A(n352), .Z(n351) );
  CIVX2 U2111 ( .A(n350), .Z(n348) );
  CIVX2 U2112 ( .A(n345), .Z(n343) );
  CIVX2 U2113 ( .A(n339), .Z(n338) );
  CIVX2 U2114 ( .A(n328), .Z(n326) );
  CIVX2 U2115 ( .A(n327), .Z(n402) );
  CIVX2 U2116 ( .A(n318), .Z(n316) );
  CIVX2 U2117 ( .A(n306), .Z(n308) );
  CIVX2 U2118 ( .A(n305), .Z(n399) );
  CIVX2 U2119 ( .A(n290), .Z(n288) );
  CIVX2 U2120 ( .A(n285), .Z(n283) );
  CIVX2 U2121 ( .A(n279), .Z(n278) );
  CIVX2 U2122 ( .A(n273), .Z(n275) );
  CIVX2 U2123 ( .A(n272), .Z(n394) );
  CIVX2 U2124 ( .A(n261), .Z(n263) );
  CIVX2 U2125 ( .A(n259), .Z(n257) );
  CIVX2 U2126 ( .A(n239), .Z(n390) );
  CIVX2 U2127 ( .A(n212), .Z(n210) );
  CIVX2 U2128 ( .A(n207), .Z(n205) );
  CIVX2 U2129 ( .A(n104), .Z(n1470) );
  CIVX2 U2130 ( .A(n109), .Z(n1469) );
  CIVX2 U2131 ( .A(n113), .Z(n1468) );
endmodule


module calc_DW_mult_uns_13 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n3, n9, n12, n15, n18, n21, n27, n30, n36, n39, n42, n44, n48, n53,
         n55, n58, n61, n63, n66, n69, n71, n74, n77, n79, n82, n85, n87, n89,
         n91, n93, n95, n97, n99, n100, n102, n104, n105, n107, n109, n110,
         n112, n113, n114, n115, n116, n120, n122, n124, n126, n128, n130,
         n132, n134, n136, n138, n140, n142, n144, n146, n148, n150, n151,
         n152, n153, n154, n155, n156, n157, n168, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n198,
         n199, n201, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n217, n218, n219, n220, n222, n225, n226, n227,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n239, n241,
         n242, n243, n244, n248, n250, n251, n252, n253, n254, n255, n259,
         n261, n262, n263, n264, n266, n270, n271, n272, n274, n276, n277,
         n278, n279, n280, n281, n282, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n297, n299, n300, n301, n302,
         n304, n307, n308, n309, n310, n312, n314, n315, n317, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n334, n336, n337, n339, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n357, n359,
         n360, n361, n362, n363, n365, n367, n368, n369, n370, n371, n373,
         n375, n376, n378, n381, n382, n383, n384, n388, n390, n391, n392,
         n394, n397, n398, n401, n402, n403, n405, n407, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1438, n1439, n1440, n1442, n1443, n1445,
         n1447, n1448, n1449, n1450, n1453, n1463, n1464, n1465, n1466, n1467,
         n1468, n1552, n1553, n1554, n1555, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739;
  assign n3 = a[1];
  assign n12 = a[3];
  assign n21 = a[5];
  assign n30 = a[7];
  assign n39 = a[9];
  assign n48 = a[11];
  assign n55 = a[13];
  assign n63 = a[15];
  assign n71 = a[17];
  assign n79 = a[19];
  assign n87 = a[21];
  assign n93 = a[23];
  assign n99 = a[25];
  assign n104 = a[27];
  assign n109 = a[29];
  assign n113 = a[31];
  assign n116 = b[0];
  assign n120 = b[1];
  assign n122 = b[2];
  assign n124 = b[3];
  assign n126 = b[4];
  assign n128 = b[5];
  assign n130 = b[6];
  assign n132 = b[7];
  assign n134 = b[8];
  assign n136 = b[9];
  assign n138 = b[10];
  assign n140 = b[11];
  assign n142 = b[12];
  assign n144 = b[13];
  assign n146 = b[14];
  assign n148 = b[15];
  assign n150 = b[16];
  assign n151 = b[17];
  assign n152 = b[18];
  assign n153 = b[19];
  assign n154 = b[20];
  assign n155 = b[21];
  assign n156 = b[22];
  assign n157 = b[23];

  CEO3X2 U403 ( .A(n429), .B(n411), .C(n427), .Z(n410) );
  CEO3X2 U404 ( .A(n431), .B(n413), .C(n412), .Z(n411) );
  CEO3X2 U405 ( .A(n415), .B(n433), .C(n414), .Z(n412) );
  CEO3X2 U406 ( .A(n437), .B(n435), .C(n416), .Z(n413) );
  CEO3X2 U407 ( .A(n439), .B(n418), .C(n417), .Z(n414) );
  CEO3X2 U408 ( .A(n422), .B(n419), .C(n441), .Z(n415) );
  CEO3X2 U411 ( .A(n424), .B(n451), .C(n447), .Z(n418) );
  CEO3X2 U412 ( .A(n1043), .B(n1071), .C(n1101), .Z(n419) );
  CEO3X2 U414 ( .A(n891), .B(n951), .C(n861), .Z(n421) );
  CEO3X2 U415 ( .A(n903), .B(n863), .C(n1017), .Z(n422) );
  CFA1X1 U418 ( .A(n430), .B(n428), .CI(n455), .CO(n425), .S(n426) );
  CFA1X1 U419 ( .A(n434), .B(n457), .CI(n432), .CO(n427), .S(n428) );
  CFA1X1 U420 ( .A(n436), .B(n459), .CI(n461), .CO(n429), .S(n430) );
  CFA1X1 U421 ( .A(n463), .B(n438), .CI(n440), .CO(n431), .S(n432) );
  CFA1X1 U422 ( .A(n467), .B(n442), .CI(n465), .CO(n433), .S(n434) );
  CFA1X1 U423 ( .A(n448), .B(n469), .CI(n446), .CO(n435), .S(n436) );
  CFA1X1 U424 ( .A(n452), .B(n444), .CI(n450), .CO(n437), .S(n438) );
  CFA1X1 U425 ( .A(n477), .B(n473), .CI(n475), .CO(n439), .S(n440) );
  CFA1X1 U426 ( .A(n1102), .B(n471), .CI(n479), .CO(n441), .S(n442) );
  CFA1X1 U427 ( .A(n868), .B(n1072), .CI(n864), .CO(n443), .S(n444) );
  CFA1X1 U428 ( .A(n918), .B(n1044), .CI(n952), .CO(n445), .S(n446) );
  CFA1X1 U429 ( .A(n874), .B(n994), .CI(n972), .CO(n447), .S(n448) );
  CFA1X1 U430 ( .A(n892), .B(n1018), .CI(n934), .CO(n449), .S(n450) );
  CFA1X1 U431 ( .A(n862), .B(n904), .CI(n882), .CO(n451), .S(n452) );
  CFA1X1 U432 ( .A(n458), .B(n456), .CI(n483), .CO(n453), .S(n454) );
  CFA1X1 U433 ( .A(n462), .B(n485), .CI(n460), .CO(n455), .S(n456) );
  CFA1X1 U434 ( .A(n464), .B(n487), .CI(n489), .CO(n457), .S(n458) );
  CFA1X1 U435 ( .A(n468), .B(n466), .CI(n491), .CO(n459), .S(n460) );
  CFA1X1 U436 ( .A(n470), .B(n493), .CI(n495), .CO(n461), .S(n462) );
  CFA1X1 U437 ( .A(n476), .B(n472), .CI(n474), .CO(n463), .S(n464) );
  CFA1X1 U438 ( .A(n501), .B(n478), .CI(n497), .CO(n465), .S(n466) );
  CFA1X1 U439 ( .A(n505), .B(n503), .CI(n499), .CO(n467), .S(n468) );
  CFA1X1 U440 ( .A(n1073), .B(n480), .CI(n1103), .CO(n469), .S(n470) );
  CFA1X1 U441 ( .A(n869), .B(n935), .CI(n893), .CO(n471), .S(n472) );
  CFA1X1 U442 ( .A(n919), .B(n1045), .CI(n865), .CO(n473), .S(n474) );
  CFA1X1 U443 ( .A(n875), .B(n995), .CI(n973), .CO(n475), .S(n476) );
  CFA1X1 U444 ( .A(n905), .B(n1019), .CI(n953), .CO(n477), .S(n478) );
  CHA1X1 U445 ( .A(n846), .B(n883), .CO(n479), .S(n480) );
  CFA1X1 U446 ( .A(n486), .B(n484), .CI(n509), .CO(n481), .S(n482) );
  CFA1X1 U447 ( .A(n513), .B(n511), .CI(n488), .CO(n483), .S(n484) );
  CFA1X1 U448 ( .A(n492), .B(n490), .CI(n515), .CO(n485), .S(n486) );
  CFA1X1 U449 ( .A(n496), .B(n494), .CI(n517), .CO(n487), .S(n488) );
  CFA1X1 U450 ( .A(n502), .B(n519), .CI(n521), .CO(n489), .S(n490) );
  CFA1X1 U451 ( .A(n504), .B(n498), .CI(n500), .CO(n491), .S(n492) );
  CFA1X1 U452 ( .A(n529), .B(n506), .CI(n523), .CO(n493), .S(n494) );
  CFA1X1 U453 ( .A(n531), .B(n527), .CI(n525), .CO(n495), .S(n496) );
  CFA1X1 U454 ( .A(n870), .B(n1104), .CI(n1074), .CO(n497), .S(n498) );
  CFA1X1 U455 ( .A(n876), .B(n996), .CI(n1653), .CO(n499), .S(n500) );
  CFA1X1 U456 ( .A(n920), .B(n1046), .CI(n954), .CO(n501), .S(n502) );
  CFA1X1 U457 ( .A(n884), .B(n1020), .CI(n974), .CO(n503), .S(n504) );
  CFA1X1 U458 ( .A(n866), .B(n894), .CI(n906), .CO(n505), .S(n506) );
  CFA1X1 U459 ( .A(n512), .B(n510), .CI(n535), .CO(n507), .S(n508) );
  CFA1X1 U460 ( .A(n516), .B(n537), .CI(n514), .CO(n509), .S(n510) );
  CFA1X1 U461 ( .A(n541), .B(n539), .CI(n518), .CO(n511), .S(n512) );
  CFA1X1 U462 ( .A(n522), .B(n520), .CI(n543), .CO(n513), .S(n514) );
  CFA1X1 U463 ( .A(n530), .B(n545), .CI(n528), .CO(n515), .S(n516) );
  CFA1X1 U464 ( .A(n547), .B(n524), .CI(n526), .CO(n517), .S(n518) );
  CFA1X1 U465 ( .A(n551), .B(n549), .CI(n553), .CO(n519), .S(n520) );
  CFA1X1 U466 ( .A(n937), .B(n555), .CI(n532), .CO(n521), .S(n522) );
  CFA1X1 U468 ( .A(n907), .B(n1075), .CI(n955), .CO(n525), .S(n526) );
  CFA1X1 U469 ( .A(n877), .B(n1021), .CI(n975), .CO(n527), .S(n528) );
  CFA1X1 U470 ( .A(n921), .B(n1047), .CI(n871), .CO(n529), .S(n530) );
  CFA1X1 U472 ( .A(n538), .B(n536), .CI(n559), .CO(n533), .S(n534) );
  CFA1X1 U473 ( .A(n563), .B(n540), .CI(n561), .CO(n535), .S(n536) );
  CFA1X1 U474 ( .A(n546), .B(n542), .CI(n544), .CO(n537), .S(n538) );
  CFA1X1 U475 ( .A(n569), .B(n565), .CI(n567), .CO(n539), .S(n540) );
  CFA1X1 U476 ( .A(n552), .B(n548), .CI(n550), .CO(n541), .S(n542) );
  CFA1X1 U477 ( .A(n571), .B(n554), .CI(n556), .CO(n543), .S(n544) );
  CFA1X1 U478 ( .A(n573), .B(n575), .CI(n577), .CO(n545), .S(n546) );
  CFA1X1 U480 ( .A(n878), .B(n1022), .CI(n998), .CO(n549), .S(n550) );
  CFA1X1 U481 ( .A(n908), .B(n1076), .CI(n956), .CO(n551), .S(n552) );
  CFA1X1 U482 ( .A(n886), .B(n1048), .CI(n976), .CO(n553), .S(n554) );
  CFA1X1 U483 ( .A(n872), .B(n922), .CI(n896), .CO(n555), .S(n556) );
  CFA1X1 U484 ( .A(n562), .B(n560), .CI(n583), .CO(n557), .S(n558) );
  CFA1X1 U485 ( .A(n587), .B(n585), .CI(n564), .CO(n559), .S(n560) );
  CFA1X1 U486 ( .A(n589), .B(n566), .CI(n568), .CO(n561), .S(n562) );
  CFA1X1 U487 ( .A(n593), .B(n570), .CI(n591), .CO(n563), .S(n564) );
  CFA1X1 U488 ( .A(n576), .B(n572), .CI(n574), .CO(n565), .S(n566) );
  CFA1X1 U489 ( .A(n597), .B(n578), .CI(n599), .CO(n567), .S(n568) );
  CFA1X1 U490 ( .A(n580), .B(n595), .CI(n601), .CO(n569), .S(n570) );
  CFA1X1 U491 ( .A(n909), .B(n1023), .CI(n957), .CO(n571), .S(n572) );
  CFA1X1 U493 ( .A(n1652), .B(n1107), .CI(n999), .CO(n575), .S(n576) );
  CHA1X1 U495 ( .A(n848), .B(n887), .CO(n579), .S(n580) );
  CFA1X1 U496 ( .A(n586), .B(n584), .CI(n605), .CO(n581), .S(n582) );
  CFA1X1 U497 ( .A(n609), .B(n588), .CI(n607), .CO(n583), .S(n584) );
  CFA1X1 U498 ( .A(n592), .B(n590), .CI(n611), .CO(n585), .S(n586) );
  CFA1X1 U499 ( .A(n598), .B(n594), .CI(n613), .CO(n587), .S(n588) );
  CFA1X1 U501 ( .A(n617), .B(n602), .CI(n621), .CO(n591), .S(n592) );
  CFA1X1 U502 ( .A(n1024), .B(n619), .CI(n623), .CO(n593), .S(n594) );
  CFA1X1 U504 ( .A(n940), .B(n1108), .CI(n978), .CO(n597), .S(n598) );
  CFA1X1 U505 ( .A(n888), .B(n1078), .CI(n1000), .CO(n599), .S(n600) );
  CFA1X1 U506 ( .A(n880), .B(n924), .CI(n898), .CO(n601), .S(n602) );
  CFA1X1 U508 ( .A(n612), .B(n629), .CI(n610), .CO(n605), .S(n606) );
  CFA1X1 U510 ( .A(n618), .B(n635), .CI(n616), .CO(n609), .S(n610) );
  CFA1X1 U511 ( .A(n639), .B(n620), .CI(n622), .CO(n611), .S(n612) );
  CFA1X1 U512 ( .A(n643), .B(n637), .CI(n641), .CO(n613), .S(n614) );
  CFA1X1 U513 ( .A(n911), .B(n1025), .CI(n624), .CO(n615), .S(n616) );
  CFA1X1 U515 ( .A(n1655), .B(n1079), .CI(n889), .CO(n619), .S(n620) );
  CFA1X1 U516 ( .A(n1001), .B(n941), .CI(n1109), .CO(n621), .S(n622) );
  CHA1X1 U517 ( .A(n899), .B(n849), .CO(n623), .S(n624) );
  CFA1X1 U518 ( .A(n630), .B(n628), .CI(n647), .CO(n625), .S(n626) );
  CFA1X1 U519 ( .A(n634), .B(n649), .CI(n632), .CO(n627), .S(n628) );
  CFA1X1 U520 ( .A(n653), .B(n651), .CI(n636), .CO(n629), .S(n630) );
  CFA1X1 U521 ( .A(n640), .B(n638), .CI(n655), .CO(n631), .S(n632) );
  CFA1X1 U522 ( .A(n659), .B(n642), .CI(n644), .CO(n633), .S(n634) );
  CFA1X1 U523 ( .A(n663), .B(n657), .CI(n661), .CO(n635), .S(n636) );
  CFA1X1 U524 ( .A(n960), .B(n1052), .CI(n1026), .CO(n637), .S(n638) );
  CFA1X1 U525 ( .A(n1654), .B(n1080), .CI(n980), .CO(n639), .S(n640) );
  CFA1X1 U526 ( .A(n912), .B(n1110), .CI(n1002), .CO(n641), .S(n642) );
  CFA1X1 U527 ( .A(n890), .B(n942), .CI(n1651), .CO(n643), .S(n644) );
  CFA1X1 U528 ( .A(n650), .B(n648), .CI(n667), .CO(n645), .S(n646) );
  CFA1X1 U529 ( .A(n654), .B(n669), .CI(n652), .CO(n647), .S(n648) );
  CFA1X1 U530 ( .A(n656), .B(n671), .CI(n673), .CO(n649), .S(n650) );
  CFA1X1 U531 ( .A(n662), .B(n658), .CI(n660), .CO(n651), .S(n652) );
  CFA1X1 U532 ( .A(n677), .B(n675), .CI(n679), .CO(n653), .S(n654) );
  CFA1X1 U533 ( .A(n901), .B(n681), .CI(n664), .CO(n655), .S(n656) );
  CFA1X1 U534 ( .A(n981), .B(n1053), .CI(n927), .CO(n657), .S(n658) );
  CFA1X1 U535 ( .A(n913), .B(n1081), .CI(n1027), .CO(n659), .S(n660) );
  CFA1X1 U536 ( .A(n961), .B(n1111), .CI(n1003), .CO(n661), .S(n662) );
  CHA1X1 U537 ( .A(n943), .B(n850), .CO(n663), .S(n664) );
  CFA1X1 U538 ( .A(n670), .B(n668), .CI(n685), .CO(n665), .S(n666) );
  CFA1X1 U539 ( .A(n674), .B(n687), .CI(n672), .CO(n667), .S(n668) );
  CFA1X1 U540 ( .A(n676), .B(n689), .CI(n691), .CO(n669), .S(n670) );
  CFA1X1 U541 ( .A(n682), .B(n678), .CI(n680), .CO(n671), .S(n672) );
  CFA1X1 U542 ( .A(n693), .B(n697), .CI(n695), .CO(n673), .S(n674) );
  CFA1X1 U543 ( .A(n1028), .B(n699), .CI(n1054), .CO(n675), .S(n676) );
  CFA1X1 U545 ( .A(n962), .B(n1112), .CI(n1004), .CO(n679), .S(n680) );
  CFA1X1 U546 ( .A(n914), .B(n944), .CI(n902), .CO(n681), .S(n682) );
  CFA1X1 U547 ( .A(n688), .B(n686), .CI(n703), .CO(n683), .S(n684) );
  CFA1X1 U548 ( .A(n692), .B(n705), .CI(n690), .CO(n685), .S(n686) );
  CFA1X1 U549 ( .A(n694), .B(n707), .CI(n709), .CO(n687), .S(n688) );
  CFA1X1 U550 ( .A(n713), .B(n696), .CI(n698), .CO(n689), .S(n690) );
  CFA1X1 U551 ( .A(n700), .B(n711), .CI(n715), .CO(n691), .S(n692) );
  CFA1X1 U552 ( .A(n929), .B(n1055), .CI(n1005), .CO(n693), .S(n694) );
  CFA1X1 U553 ( .A(n945), .B(n1083), .CI(n915), .CO(n695), .S(n696) );
  CFA1X1 U554 ( .A(n1029), .B(n1113), .CI(n983), .CO(n697), .S(n698) );
  CHA1X1 U555 ( .A(n851), .B(n963), .CO(n699), .S(n700) );
  CFA1X1 U556 ( .A(n706), .B(n704), .CI(n719), .CO(n701), .S(n702) );
  CFA1X1 U557 ( .A(n710), .B(n721), .CI(n708), .CO(n703), .S(n704) );
  CFA1X1 U558 ( .A(n712), .B(n723), .CI(n725), .CO(n705), .S(n706) );
  CFA1X1 U559 ( .A(n729), .B(n714), .CI(n716), .CO(n707), .S(n708) );
  CFA1X1 U560 ( .A(n1056), .B(n727), .CI(n731), .CO(n709), .S(n710) );
  CFA1X1 U561 ( .A(n984), .B(n1084), .CI(n1006), .CO(n711), .S(n712) );
  CFA1X1 U562 ( .A(n946), .B(n1114), .CI(n1030), .CO(n713), .S(n714) );
  CFA1X1 U563 ( .A(n916), .B(n930), .CI(n964), .CO(n715), .S(n716) );
  CFA1X1 U564 ( .A(n722), .B(n720), .CI(n735), .CO(n717), .S(n718) );
  CFA1X1 U565 ( .A(n739), .B(n737), .CI(n724), .CO(n719), .S(n720) );
  CFA1X1 U566 ( .A(n730), .B(n726), .CI(n728), .CO(n721), .S(n722) );
  CFA1X1 U567 ( .A(n745), .B(n741), .CI(n743), .CO(n723), .S(n724) );
  CFA1X1 U568 ( .A(n947), .B(n732), .CI(n1057), .CO(n725), .S(n726) );
  CFA1X1 U569 ( .A(n965), .B(n1085), .CI(n931), .CO(n727), .S(n728) );
  CFA1X1 U570 ( .A(n985), .B(n1115), .CI(n1031), .CO(n729), .S(n730) );
  CHA1X1 U571 ( .A(n852), .B(n1007), .CO(n731), .S(n732) );
  CFA1X1 U572 ( .A(n738), .B(n736), .CI(n749), .CO(n733), .S(n734) );
  CFA1X1 U573 ( .A(n753), .B(n751), .CI(n740), .CO(n735), .S(n736) );
  CFA1X1 U574 ( .A(n746), .B(n742), .CI(n744), .CO(n737), .S(n738) );
  CFA1X1 U575 ( .A(n759), .B(n755), .CI(n757), .CO(n739), .S(n740) );
  CFA1X1 U576 ( .A(n1008), .B(n1086), .CI(n1058), .CO(n741), .S(n742) );
  CFA1X1 U577 ( .A(n948), .B(n1116), .CI(n1032), .CO(n743), .S(n744) );
  CFA1X1 U578 ( .A(n932), .B(n986), .CI(n966), .CO(n745), .S(n746) );
  CFA1X1 U579 ( .A(n752), .B(n750), .CI(n763), .CO(n747), .S(n748) );
  CFA1X1 U580 ( .A(n756), .B(n754), .CI(n765), .CO(n749), .S(n750) );
  CFA1X1 U581 ( .A(n769), .B(n758), .CI(n767), .CO(n751), .S(n752) );
  CFA1X1 U582 ( .A(n967), .B(n771), .CI(n760), .CO(n753), .S(n754) );
  CFA1X1 U583 ( .A(n1009), .B(n1087), .CI(n1059), .CO(n755), .S(n756) );
  CFA1X1 U584 ( .A(n987), .B(n1117), .CI(n1033), .CO(n757), .S(n758) );
  CHA1X1 U585 ( .A(n853), .B(n949), .CO(n759), .S(n760) );
  CFA1X1 U586 ( .A(n766), .B(n764), .CI(n775), .CO(n761), .S(n762) );
  CFA1X1 U587 ( .A(n770), .B(n777), .CI(n768), .CO(n763), .S(n764) );
  CFA1X1 U588 ( .A(n779), .B(n772), .CI(n781), .CO(n765), .S(n766) );
  CFA1X1 U589 ( .A(n1034), .B(n783), .CI(n1088), .CO(n767), .S(n768) );
  CFA1X1 U590 ( .A(n1010), .B(n1118), .CI(n1060), .CO(n769), .S(n770) );
  CFA1X1 U591 ( .A(n950), .B(n968), .CI(n988), .CO(n771), .S(n772) );
  CFA1X1 U592 ( .A(n778), .B(n776), .CI(n787), .CO(n773), .S(n774) );
  CFA1X1 U593 ( .A(n782), .B(n789), .CI(n780), .CO(n775), .S(n776) );
  CFA1X1 U594 ( .A(n784), .B(n791), .CI(n793), .CO(n777), .S(n778) );
  CFA1X1 U595 ( .A(n989), .B(n1089), .CI(n969), .CO(n779), .S(n780) );
  CFA1X1 U596 ( .A(n1011), .B(n1119), .CI(n1061), .CO(n781), .S(n782) );
  CHA1X1 U597 ( .A(n854), .B(n1035), .CO(n783), .S(n784) );
  CFA1X1 U598 ( .A(n797), .B(n788), .CI(n790), .CO(n785), .S(n786) );
  CFA1X1 U599 ( .A(n794), .B(n799), .CI(n792), .CO(n787), .S(n788) );
  CFA1X1 U600 ( .A(n1062), .B(n801), .CI(n803), .CO(n789), .S(n790) );
  CFA1X1 U601 ( .A(n1036), .B(n1120), .CI(n1090), .CO(n791), .S(n792) );
  CFA1X1 U602 ( .A(n970), .B(n1012), .CI(n990), .CO(n793), .S(n794) );
  CFA1X1 U603 ( .A(n800), .B(n798), .CI(n807), .CO(n795), .S(n796) );
  CFA1X1 U604 ( .A(n811), .B(n802), .CI(n809), .CO(n797), .S(n798) );
  CFA1X1 U605 ( .A(n991), .B(n804), .CI(n1091), .CO(n799), .S(n800) );
  CFA1X1 U606 ( .A(n1013), .B(n1121), .CI(n1063), .CO(n801), .S(n802) );
  CHA1X1 U607 ( .A(n855), .B(n1037), .CO(n803), .S(n804) );
  CFA1X1 U608 ( .A(n810), .B(n808), .CI(n815), .CO(n805), .S(n806) );
  CFA1X1 U609 ( .A(n819), .B(n812), .CI(n817), .CO(n807), .S(n808) );
  CFA1X1 U610 ( .A(n1064), .B(n1122), .CI(n1092), .CO(n809), .S(n810) );
  CFA1X1 U611 ( .A(n992), .B(n1038), .CI(n1014), .CO(n811), .S(n812) );
  CFA1X1 U612 ( .A(n818), .B(n816), .CI(n823), .CO(n813), .S(n814) );
  CFA1X1 U613 ( .A(n1039), .B(n825), .CI(n820), .CO(n815), .S(n816) );
  CFA1X1 U614 ( .A(n1015), .B(n1123), .CI(n1065), .CO(n817), .S(n818) );
  CHA1X1 U615 ( .A(n856), .B(n1093), .CO(n819), .S(n820) );
  CFA1X1 U616 ( .A(n829), .B(n824), .CI(n826), .CO(n821), .S(n822) );
  CFA1X1 U617 ( .A(n1094), .B(n831), .CI(n1124), .CO(n823), .S(n824) );
  CFA1X1 U618 ( .A(n1016), .B(n1066), .CI(n1040), .CO(n825), .S(n826) );
  CFA1X1 U619 ( .A(n832), .B(n830), .CI(n835), .CO(n827), .S(n828) );
  CFA1X1 U620 ( .A(n1041), .B(n1095), .CI(n1067), .CO(n829), .S(n830) );
  CHA1X1 U621 ( .A(n857), .B(n1125), .CO(n831), .S(n832) );
  CFA1X1 U622 ( .A(n1126), .B(n836), .CI(n839), .CO(n833), .S(n834) );
  CFA1X1 U623 ( .A(n1042), .B(n1096), .CI(n1591), .CO(n835), .S(n836) );
  CFA1X1 U624 ( .A(n1069), .B(n840), .CI(n1097), .CO(n837), .S(n838) );
  CHA1X1 U625 ( .A(n858), .B(n1127), .CO(n839), .S(n840) );
  CFA1X1 U626 ( .A(n1070), .B(n1128), .CI(n1098), .CO(n841), .S(n842) );
  CHA1X1 U627 ( .A(n859), .B(n1099), .CO(n843), .S(n844) );
  COND2X1 U628 ( .A(n115), .B(n1463), .C(n114), .D(n1134), .Z(n845) );
  COND2X1 U629 ( .A(n1132), .B(n114), .C(n115), .D(n1133), .Z(n861) );
  CND2IX1 U633 ( .B(n1691), .A(n113), .Z(n1134) );
  COND2X1 U634 ( .A(n112), .B(n1464), .C(n110), .D(n1139), .Z(n846) );
  COND2X1 U635 ( .A(n1135), .B(n110), .C(n1136), .D(n112), .Z(n863) );
  COND2X1 U636 ( .A(n1137), .B(n112), .C(n110), .D(n1136), .Z(n864) );
  COND2X1 U637 ( .A(n1137), .B(n110), .C(n112), .D(n1138), .Z(n865) );
  COND2X1 U644 ( .A(n107), .B(n1465), .C(n105), .D(n1146), .Z(n847) );
  COND2X1 U645 ( .A(n1140), .B(n105), .C(n1141), .D(n107), .Z(n867) );
  COND2X1 U646 ( .A(n1142), .B(n107), .C(n105), .D(n1141), .Z(n868) );
  COND2X1 U647 ( .A(n1142), .B(n105), .C(n1143), .D(n107), .Z(n869) );
  COND2X1 U648 ( .A(n1144), .B(n107), .C(n105), .D(n1143), .Z(n870) );
  CND2IX1 U657 ( .B(n1691), .A(n104), .Z(n1146) );
  COND2X1 U658 ( .A(n102), .B(n1466), .C(n100), .D(n1155), .Z(n848) );
  COND2X1 U660 ( .A(n1149), .B(n102), .C(n100), .D(n1148), .Z(n874) );
  COND2X1 U661 ( .A(n1149), .B(n100), .C(n1150), .D(n102), .Z(n875) );
  COND2X1 U662 ( .A(n1151), .B(n102), .C(n100), .D(n1150), .Z(n876) );
  COND2X1 U663 ( .A(n1151), .B(n100), .C(n1152), .D(n102), .Z(n877) );
  COND2X1 U664 ( .A(n1153), .B(n102), .C(n100), .D(n1152), .Z(n878) );
  COND2X1 U676 ( .A(n97), .B(n1467), .C(n95), .D(n1166), .Z(n849) );
  COND2X1 U680 ( .A(n1160), .B(n97), .C(n1159), .D(n95), .Z(n884) );
  COND2X1 U683 ( .A(n1162), .B(n95), .C(n1163), .D(n97), .Z(n887) );
  COND2X1 U684 ( .A(n1164), .B(n97), .C(n1163), .D(n95), .Z(n888) );
  COND2X1 U685 ( .A(n1164), .B(n95), .C(n97), .D(n1165), .Z(n889) );
  CND2IX1 U697 ( .B(n1691), .A(n1688), .Z(n1166) );
  COND2X1 U727 ( .A(n85), .B(n1183), .C(n1657), .D(n1182), .Z(n905) );
  COND2X1 U729 ( .A(n85), .B(n1185), .C(n1657), .D(n1184), .Z(n907) );
  COND2X1 U730 ( .A(n85), .B(n1186), .C(n1185), .D(n1657), .Z(n908) );
  COND2X1 U731 ( .A(n85), .B(n1187), .C(n1657), .D(n1186), .Z(n909) );
  COND2X1 U732 ( .A(n1188), .B(n85), .C(n1187), .D(n1657), .Z(n910) );
  COND2X1 U734 ( .A(n1190), .B(n85), .C(n1189), .D(n1657), .Z(n912) );
  COND2X1 U737 ( .A(n1193), .B(n85), .C(n1657), .D(n1192), .Z(n915) );
  COND2X1 U797 ( .A(n69), .B(n1221), .C(n66), .D(n1220), .Z(n941) );
  COND2X1 U799 ( .A(n69), .B(n1223), .C(n66), .D(n1222), .Z(n943) );
  COND2X1 U800 ( .A(n69), .B(n1224), .C(n1223), .D(n66), .Z(n944) );
  COND2X1 U801 ( .A(n69), .B(n1225), .C(n66), .D(n1224), .Z(n945) );
  COND2X1 U802 ( .A(n69), .B(n1226), .C(n1225), .D(n66), .Z(n946) );
  COND2X1 U804 ( .A(n69), .B(n1228), .C(n1227), .D(n66), .Z(n948) );
  COND2X1 U829 ( .A(n61), .B(n1234), .C(n58), .D(n1233), .Z(n953) );
  COND2X1 U830 ( .A(n61), .B(n1235), .C(n1234), .D(n58), .Z(n954) );
  COND2X1 U831 ( .A(n61), .B(n1236), .C(n58), .D(n1235), .Z(n955) );
  COND2X1 U832 ( .A(n61), .B(n1237), .C(n1236), .D(n58), .Z(n956) );
  COND2X1 U833 ( .A(n61), .B(n1238), .C(n58), .D(n1237), .Z(n957) );
  COND2X1 U834 ( .A(n61), .B(n1239), .C(n1238), .D(n58), .Z(n958) );
  COND2X1 U835 ( .A(n61), .B(n1240), .C(n58), .D(n1239), .Z(n959) );
  COND2X1 U836 ( .A(n61), .B(n1241), .C(n1240), .D(n58), .Z(n960) );
  COND2X1 U837 ( .A(n61), .B(n1242), .C(n58), .D(n1241), .Z(n961) );
  COND2X1 U838 ( .A(n61), .B(n1243), .C(n1242), .D(n58), .Z(n962) );
  COND2X1 U839 ( .A(n61), .B(n1244), .C(n58), .D(n1243), .Z(n963) );
  COND2X1 U840 ( .A(n61), .B(n1245), .C(n1244), .D(n58), .Z(n964) );
  COND2X1 U841 ( .A(n61), .B(n1246), .C(n58), .D(n1245), .Z(n965) );
  COND2X1 U842 ( .A(n61), .B(n1247), .C(n1246), .D(n58), .Z(n966) );
  COND2X1 U844 ( .A(n61), .B(n1249), .C(n1248), .D(n58), .Z(n968) );
  COND2X1 U845 ( .A(n61), .B(n1250), .C(n58), .D(n1249), .Z(n969) );
  COND2X1 U871 ( .A(n53), .B(n1255), .C(n1254), .D(n1624), .Z(n973) );
  COND2X1 U872 ( .A(n53), .B(n1256), .C(n1255), .D(n1624), .Z(n974) );
  COND2X1 U873 ( .A(n53), .B(n1257), .C(n1624), .D(n1256), .Z(n975) );
  COND2X1 U874 ( .A(n53), .B(n1258), .C(n1257), .D(n1624), .Z(n976) );
  COND2X1 U876 ( .A(n53), .B(n1260), .C(n1259), .D(n1624), .Z(n978) );
  COND2X1 U877 ( .A(n53), .B(n1261), .C(n1624), .D(n1260), .Z(n979) );
  COND2X1 U878 ( .A(n53), .B(n1262), .C(n1261), .D(n1624), .Z(n980) );
  COND2X1 U879 ( .A(n53), .B(n1263), .C(n1624), .D(n1262), .Z(n981) );
  COND2X1 U880 ( .A(n53), .B(n1264), .C(n1263), .D(n1624), .Z(n982) );
  COND2X1 U881 ( .A(n53), .B(n1265), .C(n1624), .D(n1264), .Z(n983) );
  COND2X1 U882 ( .A(n53), .B(n1266), .C(n1265), .D(n1624), .Z(n984) );
  COND2X1 U884 ( .A(n53), .B(n1268), .C(n1267), .D(n1624), .Z(n986) );
  COND2X1 U885 ( .A(n53), .B(n1269), .C(n1624), .D(n1268), .Z(n987) );
  COND2X1 U886 ( .A(n53), .B(n1270), .C(n1269), .D(n1624), .Z(n988) );
  COND2X1 U887 ( .A(n53), .B(n1271), .C(n1624), .D(n1270), .Z(n989) );
  COND2X1 U888 ( .A(n53), .B(n1272), .C(n1271), .D(n1624), .Z(n990) );
  CND2IX1 U913 ( .B(n1691), .A(n1722), .Z(n1274) );
  COND2X1 U914 ( .A(n44), .B(n1718), .C(n1299), .D(n42), .Z(n856) );
  COND2X1 U915 ( .A(n1555), .B(n1276), .C(n1275), .D(n42), .Z(n993) );
  COND2X1 U916 ( .A(n1555), .B(n1277), .C(n1276), .D(n42), .Z(n994) );
  COND2X1 U917 ( .A(n1555), .B(n1278), .C(n1277), .D(n42), .Z(n995) );
  COND2X1 U920 ( .A(n44), .B(n1281), .C(n1280), .D(n42), .Z(n998) );
  COND2X1 U922 ( .A(n44), .B(n1283), .C(n1282), .D(n42), .Z(n1000) );
  COND2X1 U923 ( .A(n44), .B(n1284), .C(n1283), .D(n42), .Z(n1001) );
  COND2X1 U924 ( .A(n44), .B(n1285), .C(n1284), .D(n42), .Z(n1002) );
  COND2X1 U925 ( .A(n44), .B(n1286), .C(n42), .D(n1285), .Z(n1003) );
  COND2X1 U926 ( .A(n44), .B(n1287), .C(n1286), .D(n42), .Z(n1004) );
  COND2X1 U928 ( .A(n1555), .B(n1289), .C(n1288), .D(n42), .Z(n1006) );
  COND2X1 U929 ( .A(n44), .B(n1290), .C(n42), .D(n1289), .Z(n1007) );
  COND2X1 U930 ( .A(n44), .B(n1291), .C(n1290), .D(n42), .Z(n1008) );
  COND2X1 U931 ( .A(n44), .B(n1292), .C(n42), .D(n1291), .Z(n1009) );
  COND2X1 U933 ( .A(n44), .B(n1294), .C(n42), .D(n1293), .Z(n1011) );
  COND2X1 U934 ( .A(n1555), .B(n1295), .C(n1294), .D(n42), .Z(n1012) );
  COND2X1 U935 ( .A(n44), .B(n1296), .C(n42), .D(n1295), .Z(n1013) );
  COND2X1 U936 ( .A(n44), .B(n1297), .C(n1296), .D(n42), .Z(n1014) );
  COND2X1 U937 ( .A(n44), .B(n1298), .C(n42), .D(n1297), .Z(n1015) );
  COND2X1 U966 ( .A(n36), .B(n1302), .C(n1301), .D(n1621), .Z(n1018) );
  COND2X1 U967 ( .A(n36), .B(n1303), .C(n1302), .D(n1621), .Z(n1019) );
  COND2X1 U968 ( .A(n36), .B(n1304), .C(n1303), .D(n1621), .Z(n1020) );
  COND2X1 U969 ( .A(n36), .B(n1305), .C(n1304), .D(n1621), .Z(n1021) );
  COND2X1 U970 ( .A(n36), .B(n1306), .C(n1305), .D(n1621), .Z(n1022) );
  COND2X1 U971 ( .A(n36), .B(n1307), .C(n1306), .D(n1621), .Z(n1023) );
  COND2X1 U972 ( .A(n36), .B(n1308), .C(n1307), .D(n1621), .Z(n1024) );
  COND2X1 U974 ( .A(n36), .B(n1310), .C(n1309), .D(n1621), .Z(n1026) );
  COND2X1 U976 ( .A(n36), .B(n1312), .C(n1311), .D(n1621), .Z(n1028) );
  COND2X1 U978 ( .A(n36), .B(n1314), .C(n1313), .D(n1621), .Z(n1030) );
  COND2X1 U980 ( .A(n36), .B(n1316), .C(n1315), .D(n1621), .Z(n1032) );
  COND2X1 U981 ( .A(n36), .B(n1317), .C(n1621), .D(n1316), .Z(n1033) );
  COND2X1 U982 ( .A(n36), .B(n1318), .C(n1317), .D(n1621), .Z(n1034) );
  COND2X1 U984 ( .A(n36), .B(n1320), .C(n1319), .D(n1621), .Z(n1036) );
  COND2X1 U985 ( .A(n36), .B(n1321), .C(n1621), .D(n1320), .Z(n1037) );
  COND2X1 U987 ( .A(n36), .B(n1323), .C(n1621), .D(n1322), .Z(n1039) );
  COND2X1 U988 ( .A(n36), .B(n1324), .C(n1323), .D(n1621), .Z(n1040) );
  CND2IX1 U1017 ( .B(n1691), .A(n1709), .Z(n1326) );
  COND2X1 U1026 ( .A(n27), .B(n1335), .C(n1334), .D(n1623), .Z(n1050) );
  COND2X1 U1028 ( .A(n27), .B(n1337), .C(n1336), .D(n1623), .Z(n1052) );
  COND2X1 U1030 ( .A(n27), .B(n1339), .C(n1338), .D(n1623), .Z(n1054) );
  COND2X1 U1033 ( .A(n27), .B(n1342), .C(n1341), .D(n1623), .Z(n1057) );
  COND2X1 U1034 ( .A(n27), .B(n1343), .C(n1342), .D(n1623), .Z(n1058) );
  COND2X1 U1035 ( .A(n27), .B(n1344), .C(n1343), .D(n1623), .Z(n1059) );
  COND2X1 U1037 ( .A(n27), .B(n1346), .C(n1623), .D(n1345), .Z(n1061) );
  COND2X1 U1039 ( .A(n27), .B(n1348), .C(n1623), .D(n1347), .Z(n1063) );
  COND2X1 U1040 ( .A(n27), .B(n1349), .C(n1348), .D(n1623), .Z(n1064) );
  COND2X1 U1041 ( .A(n27), .B(n1350), .C(n1623), .D(n1349), .Z(n1065) );
  COND2X1 U1077 ( .A(n18), .B(n1357), .C(n1356), .D(n15), .Z(n1071) );
  COND2X1 U1078 ( .A(n18), .B(n1358), .C(n1357), .D(n15), .Z(n1072) );
  COND2X1 U1079 ( .A(n18), .B(n1359), .C(n1358), .D(n15), .Z(n1073) );
  COND2X1 U1080 ( .A(n18), .B(n1360), .C(n1359), .D(n15), .Z(n1074) );
  COND2X1 U1081 ( .A(n18), .B(n1361), .C(n1360), .D(n15), .Z(n1075) );
  COND2X1 U1082 ( .A(n18), .B(n1362), .C(n1361), .D(n15), .Z(n1076) );
  COND2X1 U1084 ( .A(n18), .B(n1364), .C(n1363), .D(n15), .Z(n1078) );
  COND2X1 U1085 ( .A(n18), .B(n1365), .C(n1364), .D(n15), .Z(n1079) );
  COND2X1 U1089 ( .A(n18), .B(n1369), .C(n1368), .D(n15), .Z(n1083) );
  COND2X1 U1090 ( .A(n18), .B(n1370), .C(n1369), .D(n15), .Z(n1084) );
  COND2X1 U1091 ( .A(n18), .B(n1371), .C(n1370), .D(n15), .Z(n1085) );
  COND2X1 U1092 ( .A(n18), .B(n1372), .C(n1371), .D(n15), .Z(n1086) );
  COND2X1 U1093 ( .A(n18), .B(n1373), .C(n1372), .D(n15), .Z(n1087) );
  COND2X1 U1094 ( .A(n18), .B(n1374), .C(n1373), .D(n15), .Z(n1088) );
  COND2X1 U1095 ( .A(n18), .B(n1375), .C(n1374), .D(n15), .Z(n1089) );
  COND2X1 U1096 ( .A(n18), .B(n1376), .C(n1375), .D(n15), .Z(n1090) );
  COND2X1 U1097 ( .A(n18), .B(n1377), .C(n15), .D(n1376), .Z(n1091) );
  COND2X1 U1098 ( .A(n18), .B(n1378), .C(n1377), .D(n15), .Z(n1092) );
  COND2X1 U1099 ( .A(n18), .B(n1379), .C(n15), .D(n1378), .Z(n1093) );
  COND2X1 U1100 ( .A(n18), .B(n1380), .C(n1379), .D(n15), .Z(n1094) );
  COND2X1 U1101 ( .A(n18), .B(n1381), .C(n15), .D(n1380), .Z(n1095) );
  COND2X1 U1102 ( .A(n18), .B(n1382), .C(n1381), .D(n15), .Z(n1096) );
  COND2X1 U1103 ( .A(n18), .B(n1383), .C(n15), .D(n1382), .Z(n1097) );
  COND2X1 U1104 ( .A(n18), .B(n1384), .C(n1383), .D(n15), .Z(n1098) );
  COND2X1 U1105 ( .A(n18), .B(n1385), .C(n15), .D(n1384), .Z(n1099) );
  COND2X1 U1138 ( .A(n1561), .B(n1599), .C(n1696), .D(n1419), .Z(n860) );
  COND2X1 U1145 ( .A(n1675), .B(n1394), .C(n1696), .D(n1393), .Z(n1107) );
  COND2X1 U1147 ( .A(n1675), .B(n1396), .C(n1696), .D(n1395), .Z(n1109) );
  COND2X1 U1149 ( .A(n1561), .B(n1398), .C(n1696), .D(n1397), .Z(n1111) );
  COND2X1 U1150 ( .A(n1675), .B(n1399), .C(n1696), .D(n1398), .Z(n1112) );
  COND2X1 U1151 ( .A(n1561), .B(n1400), .C(n1696), .D(n1399), .Z(n1113) );
  COND2X1 U1152 ( .A(n1561), .B(n1401), .C(n1696), .D(n1400), .Z(n1114) );
  COND2X1 U1153 ( .A(n1561), .B(n1402), .C(n1696), .D(n1401), .Z(n1115) );
  COND2X1 U1154 ( .A(n1561), .B(n1403), .C(n1696), .D(n1402), .Z(n1116) );
  COND2X1 U1155 ( .A(n1561), .B(n1404), .C(n1696), .D(n1403), .Z(n1117) );
  COND2X1 U1156 ( .A(n1561), .B(n1405), .C(n1696), .D(n1404), .Z(n1118) );
  COND2X1 U1157 ( .A(n1561), .B(n1406), .C(n1696), .D(n1405), .Z(n1119) );
  COND2X1 U1158 ( .A(n1561), .B(n1407), .C(n1696), .D(n1406), .Z(n1120) );
  COND2X1 U1159 ( .A(n1561), .B(n1408), .C(n1696), .D(n1407), .Z(n1121) );
  COND2X1 U1162 ( .A(n1561), .B(n1411), .C(n1696), .D(n1410), .Z(n1124) );
  COND2X1 U1163 ( .A(n1561), .B(n1412), .C(n1696), .D(n1411), .Z(n1125) );
  COND2X1 U1164 ( .A(n1561), .B(n1413), .C(n1696), .D(n1412), .Z(n1126) );
  COND2X1 U1165 ( .A(n1561), .B(n1414), .C(n1696), .D(n1413), .Z(n1127) );
  COND2X1 U1167 ( .A(n1561), .B(n1416), .C(n1696), .D(n1415), .Z(n1129) );
  COND2X1 U1168 ( .A(n1561), .B(n1417), .C(n1696), .D(n1416), .Z(n1130) );
  COND2X1 U1169 ( .A(n1561), .B(n1418), .C(n1696), .D(n1417), .Z(n1131) );
  CND2IX1 U1203 ( .B(n1691), .A(n1589), .Z(n1419) );
  COND2X1 U1276 ( .A(n1192), .B(n85), .C(n1191), .D(n82), .Z(n914) );
  CND2IX4 U1277 ( .B(n1619), .A(n82), .Z(n85) );
  CND2X1 U1278 ( .A(n1578), .B(n1579), .Z(n1192) );
  CFA1X2 U1279 ( .A(n959), .B(n1051), .CI(n979), .CO(n617), .S(n618) );
  CANR1X2 U1280 ( .A(n1635), .B(n279), .C(n274), .Z(n1552) );
  CIVX3 U1281 ( .A(n1614), .Z(n1628) );
  CNIVX2 U1282 ( .A(n140), .Z(n1684) );
  CNIVX2 U1283 ( .A(n936), .Z(n1653) );
  COND2XL U1284 ( .A(n1147), .B(n100), .C(n1148), .D(n102), .Z(n873) );
  CHA1X1 U1285 ( .A(n847), .B(n885), .CO(n531), .S(n532) );
  CANR1XL U1286 ( .A(n1635), .B(n279), .C(n274), .Z(n272) );
  COND2XL U1287 ( .A(n61), .B(n1248), .C(n58), .D(n1247), .Z(n967) );
  COR2X1 U1288 ( .A(n1202), .B(n1557), .Z(n1572) );
  CENX2 U1289 ( .A(n1687), .B(n1676), .Z(n1176) );
  CIVXL U1290 ( .A(n288), .Z(n287) );
  CND2X4 U1291 ( .A(n74), .B(n1445), .Z(n77) );
  CEOX1 U1292 ( .A(a[10]), .B(n1721), .Z(n1448) );
  CENX1 U1293 ( .A(n1682), .B(n1707), .Z(n1345) );
  CNIVX2 U1294 ( .A(n136), .Z(n1682) );
  CND2X4 U1295 ( .A(n1449), .B(n42), .Z(n44) );
  CENXL U1296 ( .A(n153), .B(n1724), .Z(n1231) );
  CENXL U1297 ( .A(n1691), .B(n1724), .Z(n1250) );
  CENXL U1298 ( .A(n1682), .B(n1724), .Z(n1241) );
  CENXL U1299 ( .A(n1694), .B(n1724), .Z(n1247) );
  CENXL U1300 ( .A(n1686), .B(n1724), .Z(n1235) );
  CENXL U1301 ( .A(n1724), .B(n1676), .Z(n1248) );
  CENXL U1302 ( .A(n1724), .B(n150), .Z(n1234) );
  CENXL U1303 ( .A(n151), .B(n1724), .Z(n1233) );
  CENXL U1304 ( .A(n1678), .B(n1724), .Z(n1245) );
  CENXL U1305 ( .A(n1724), .B(n1677), .Z(n1246) );
  CENXL U1306 ( .A(n1680), .B(n1724), .Z(n1243) );
  CENXL U1307 ( .A(n1684), .B(n1724), .Z(n1239) );
  CENXL U1308 ( .A(n1724), .B(n1679), .Z(n1244) );
  CENXL U1309 ( .A(n1724), .B(n146), .Z(n1236) );
  CENXL U1310 ( .A(n1724), .B(n142), .Z(n1238) );
  CENXL U1311 ( .A(n1685), .B(n1724), .Z(n1237) );
  CENXL U1312 ( .A(n1724), .B(n1683), .Z(n1240) );
  CENXL U1313 ( .A(n1724), .B(n1681), .Z(n1242) );
  CENXL U1314 ( .A(n1701), .B(n155), .Z(n1364) );
  CENXL U1315 ( .A(n1697), .B(n155), .Z(n1397) );
  CENXL U1316 ( .A(n1690), .B(n1687), .Z(n1178) );
  CENXL U1317 ( .A(n1690), .B(n104), .Z(n1145) );
  CNIVX2 U1318 ( .A(n116), .Z(n1690) );
  CENXL U1319 ( .A(n1692), .B(n1704), .Z(n1384) );
  CENXL U1320 ( .A(n1692), .B(n1590), .Z(n1417) );
  CENXL U1321 ( .A(n1692), .B(n1722), .Z(n1272) );
  CENXL U1322 ( .A(n1692), .B(n1717), .Z(n1297) );
  CENXL U1323 ( .A(n1692), .B(n1724), .Z(n1249) );
  CENXL U1324 ( .A(n1692), .B(n1727), .Z(n1228) );
  CENXL U1325 ( .A(n1702), .B(b[29]), .Z(n1356) );
  CNIVX2 U1326 ( .A(n138), .Z(n1683) );
  CIVX3 U1327 ( .A(n1739), .Z(n1735) );
  COND2X1 U1328 ( .A(n1144), .B(n105), .C(n107), .D(n1145), .Z(n871) );
  CNIVX3 U1329 ( .A(n124), .Z(n1694) );
  CNIVX16 U1330 ( .A(n93), .Z(n1688) );
  CENX1 U1331 ( .A(n1687), .B(n1683), .Z(n1168) );
  CNIVX1 U1332 ( .A(n9), .Z(n1675) );
  CAN2X1 U1333 ( .A(n1626), .B(n1627), .Z(n253) );
  CENX1 U1334 ( .A(n1676), .B(n1689), .Z(n1152) );
  CENX1 U1335 ( .A(n1684), .B(n1710), .Z(n1314) );
  CENX1 U1336 ( .A(n1692), .B(n1732), .Z(n1209) );
  CENX1 U1337 ( .A(n1694), .B(n1727), .Z(n1226) );
  CENX1 U1338 ( .A(n1709), .B(n146), .Z(n1311) );
  CENX1 U1339 ( .A(n1692), .B(n1688), .Z(n1164) );
  CIVX2 U1340 ( .A(n48), .Z(n1723) );
  CENX1 U1341 ( .A(n1694), .B(n1689), .Z(n1151) );
  CENX1 U1342 ( .A(n1710), .B(n155), .Z(n1304) );
  CENX1 U1343 ( .A(n1680), .B(n1687), .Z(n1171) );
  CENX1 U1344 ( .A(n1677), .B(n1689), .Z(n1150) );
  CENX1 U1345 ( .A(n1687), .B(n1681), .Z(n1170) );
  CENX1 U1346 ( .A(n1692), .B(n1712), .Z(n1324) );
  CIVX3 U1347 ( .A(n1656), .Z(n42) );
  CENX1 U1348 ( .A(n1717), .B(n155), .Z(n1277) );
  CENX1 U1349 ( .A(a[24]), .B(n1689), .Z(n1625) );
  CENX1 U1350 ( .A(n1697), .B(b[29]), .Z(n1389) );
  CND2IX2 U1351 ( .B(n1649), .A(n66), .Z(n69) );
  CND2X1 U1352 ( .A(n1582), .B(n1583), .Z(n1649) );
  CND2X1 U1353 ( .A(n1580), .B(n1581), .Z(n1583) );
  CENX1 U1354 ( .A(n1682), .B(n1687), .Z(n1169) );
  CNIVX1 U1355 ( .A(n1068), .Z(n1591) );
  CND2X1 U1356 ( .A(n1453), .B(n1696), .Z(n9) );
  CENX1 U1357 ( .A(n600), .B(n615), .Z(n1644) );
  CENX1 U1358 ( .A(n1684), .B(n1687), .Z(n1167) );
  CIVX4 U1359 ( .A(n1660), .Z(n15) );
  CENX1 U1360 ( .A(n1690), .B(n1708), .Z(n1354) );
  CNIVX3 U1361 ( .A(n9), .Z(n1561) );
  CNIVX2 U1362 ( .A(n116), .Z(n1691) );
  CENX1 U1363 ( .A(n293), .B(n179), .Z(product[18]) );
  CENX1 U1364 ( .A(n251), .B(n173), .Z(product[24]) );
  CIVDX1 U1365 ( .A(n21), .Z0(n1553), .Z1(n1554) );
  CIVX2 U1366 ( .A(n1705), .Z(n1702) );
  CIVX2 U1367 ( .A(n1719), .Z(n1716) );
  CIVX2 U1368 ( .A(n30), .Z(n1713) );
  CIVX2 U1369 ( .A(a[0]), .Z(n1696) );
  CNIVX1 U1370 ( .A(n44), .Z(n1555) );
  COND2X1 U1371 ( .A(n1162), .B(n97), .C(n1161), .D(n95), .Z(n886) );
  CAN2X1 U1372 ( .A(n1618), .B(n378), .Z(product[1]) );
  CENX1 U1373 ( .A(n1687), .B(n1679), .Z(n1172) );
  CND2X1 U1374 ( .A(n508), .B(n533), .Z(n226) );
  CNIVX2 U1375 ( .A(n925), .Z(n1655) );
  COND2X1 U1376 ( .A(n1209), .B(n77), .C(n1208), .D(n1557), .Z(n930) );
  COND1X1 U1377 ( .A(n286), .B(n280), .C(n281), .Z(n279) );
  CIVX1 U1378 ( .A(n280), .Z(n390) );
  CFA1X1 U1379 ( .A(n938), .B(n579), .CI(n1106), .CO(n547), .S(n548) );
  CND2XL U1380 ( .A(n1632), .B(n261), .Z(n174) );
  CAN2XL U1381 ( .A(n382), .B(n217), .Z(n1616) );
  COND2X1 U1382 ( .A(n18), .B(n1366), .C(n1365), .D(n15), .Z(n1080) );
  COND2XL U1383 ( .A(n61), .B(n1232), .C(n58), .D(n1231), .Z(n951) );
  COND2XL U1384 ( .A(n61), .B(n1233), .C(n1232), .D(n58), .Z(n952) );
  CND2IXL U1385 ( .B(n1691), .A(n1687), .Z(n1179) );
  CENX2 U1386 ( .A(n1694), .B(n1687), .Z(n1175) );
  CEOX4 U1387 ( .A(a[20]), .B(n1687), .Z(n1443) );
  CND2X1 U1388 ( .A(n1574), .B(n1575), .Z(n1449) );
  CND2X1 U1389 ( .A(n1573), .B(n1716), .Z(n1575) );
  COND2XL U1390 ( .A(n53), .B(n1253), .C(n1252), .D(n1624), .Z(n971) );
  COND2XL U1391 ( .A(n53), .B(n1254), .C(n1253), .D(n1624), .Z(n972) );
  COND2XL U1392 ( .A(n53), .B(n1273), .C(n1624), .D(n1272), .Z(n991) );
  COND2XL U1393 ( .A(n53), .B(n1723), .C(n1274), .D(n1624), .Z(n855) );
  COND2X1 U1394 ( .A(n1561), .B(n1397), .C(n1696), .D(n1396), .Z(n1110) );
  CND2X2 U1395 ( .A(n1630), .B(n1631), .Z(n1557) );
  CND2X2 U1396 ( .A(n1630), .B(n1631), .Z(n74) );
  CNIVXL U1397 ( .A(n923), .Z(n1558) );
  CENX1 U1398 ( .A(n1559), .B(n879), .Z(n578) );
  CENX1 U1399 ( .A(n1077), .B(n923), .Z(n1559) );
  CIVX3 U1400 ( .A(n1734), .Z(n1729) );
  CND2IXL U1401 ( .B(n1691), .A(n1729), .Z(n1211) );
  CENXL U1402 ( .A(n1678), .B(n1726), .Z(n1224) );
  CIVX4 U1403 ( .A(n1728), .Z(n1726) );
  CNR2X2 U1404 ( .A(n702), .B(n717), .Z(n291) );
  CNR2IX1 U1405 ( .B(n1691), .A(n114), .Z(n862) );
  COND2XL U1406 ( .A(n77), .B(n1197), .C(n1196), .D(n1557), .Z(n918) );
  COND2XL U1407 ( .A(n77), .B(n1210), .C(n1557), .D(n1209), .Z(n931) );
  COND2XL U1408 ( .A(n77), .B(n1202), .C(n1557), .D(n1201), .Z(n923) );
  CIVX3 U1409 ( .A(n63), .Z(n1728) );
  CENX2 U1410 ( .A(n1729), .B(a[18]), .Z(n82) );
  CND2X4 U1411 ( .A(n95), .B(n1442), .Z(n97) );
  CEOX4 U1412 ( .A(a[22]), .B(n1688), .Z(n1442) );
  COND2XL U1413 ( .A(n69), .B(n1227), .C(n66), .D(n1226), .Z(n947) );
  COND2XL U1414 ( .A(n69), .B(n1222), .C(n1221), .D(n66), .Z(n942) );
  COND1X1 U1415 ( .A(n291), .B(n295), .C(n292), .Z(n290) );
  CENX2 U1416 ( .A(n1735), .B(a[20]), .Z(n89) );
  CND2X2 U1417 ( .A(n1707), .B(a[6]), .Z(n1611) );
  CANR1XL U1418 ( .A(n220), .B(n207), .C(n208), .Z(n1560) );
  CEO3XL U1419 ( .A(n631), .B(n614), .C(n633), .Z(n608) );
  CENXL U1420 ( .A(n1716), .B(n150), .Z(n1282) );
  CENXL U1421 ( .A(n1716), .B(n146), .Z(n1284) );
  CENXL U1422 ( .A(n1716), .B(n142), .Z(n1286) );
  COND2X1 U1423 ( .A(n44), .B(n1282), .C(n1281), .D(n42), .Z(n999) );
  CIVX1 U1424 ( .A(n1713), .Z(n1709) );
  COND2XL U1425 ( .A(n36), .B(n1713), .C(n1326), .D(n1621), .Z(n857) );
  CND2X1 U1426 ( .A(n1440), .B(n105), .Z(n107) );
  CEOX1 U1427 ( .A(a[26]), .B(n104), .Z(n1440) );
  CEOX1 U1428 ( .A(a[0]), .B(n1598), .Z(n1453) );
  CENX2 U1429 ( .A(n1599), .B(a[2]), .Z(n1660) );
  CNR2IX1 U1430 ( .B(n1691), .A(n100), .Z(n880) );
  CANR1X2 U1431 ( .A(n248), .B(n1640), .C(n239), .Z(n237) );
  COND2X1 U1432 ( .A(n36), .B(n1315), .C(n1621), .D(n1314), .Z(n1031) );
  CENX4 U1433 ( .A(n1687), .B(a[22]), .Z(n95) );
  CIVXL U1434 ( .A(n321), .Z(n320) );
  CND2X2 U1435 ( .A(n1628), .B(n1629), .Z(n1631) );
  CEOX1 U1436 ( .A(n928), .B(n982), .Z(n1562) );
  CEOX1 U1437 ( .A(n1562), .B(n1082), .Z(n678) );
  CND2X1 U1438 ( .A(n1082), .B(n982), .Z(n1563) );
  CND2XL U1439 ( .A(n928), .B(n1082), .Z(n1564) );
  CND2XL U1440 ( .A(n982), .B(n928), .Z(n1565) );
  CND3XL U1441 ( .A(n1563), .B(n1564), .C(n1565), .Z(n677) );
  COND2XL U1442 ( .A(n1207), .B(n77), .C(n1206), .D(n1557), .Z(n928) );
  CND2XL U1443 ( .A(n1692), .B(n1738), .Z(n1578) );
  CENXL U1444 ( .A(n1692), .B(n1554), .Z(n1353) );
  CENXL U1445 ( .A(n1692), .B(n1687), .Z(n1177) );
  CANR1XL U1446 ( .A(n234), .B(n270), .C(n235), .Z(n1592) );
  COND1X1 U1447 ( .A(n214), .B(n222), .C(n217), .Z(n213) );
  CND2XL U1448 ( .A(n1638), .B(n1637), .Z(n309) );
  CIVX4 U1449 ( .A(n1723), .Z(n1721) );
  CND2X2 U1450 ( .A(a[8]), .B(n1718), .Z(n1574) );
  CNR2X2 U1451 ( .A(n482), .B(n507), .Z(n214) );
  COND2X1 U1452 ( .A(n69), .B(n1220), .C(n1219), .D(n66), .Z(n940) );
  CENXL U1453 ( .A(n1684), .B(n1707), .Z(n1343) );
  CENXL U1454 ( .A(n1707), .B(n156), .Z(n1332) );
  CENXL U1455 ( .A(n1707), .B(n146), .Z(n1340) );
  CENXL U1456 ( .A(n1707), .B(n152), .Z(n1336) );
  CENXL U1457 ( .A(n1707), .B(n1686), .Z(n1339) );
  CENXL U1458 ( .A(n1707), .B(n154), .Z(n1334) );
  CENXL U1459 ( .A(n1707), .B(n153), .Z(n1335) );
  CENXL U1460 ( .A(n1680), .B(n1707), .Z(n1347) );
  CENX1 U1461 ( .A(a[4]), .B(n1707), .Z(n1622) );
  COND1X1 U1462 ( .A(n288), .B(n271), .C(n1552), .Z(n270) );
  CANR1X1 U1463 ( .A(n317), .B(n1638), .C(n312), .Z(n310) );
  COR2XL U1464 ( .A(n748), .B(n761), .Z(n1638) );
  CEOX1 U1465 ( .A(a[6]), .B(n30), .Z(n1450) );
  CNIVX2 U1466 ( .A(n897), .Z(n1652) );
  CNR2X1 U1467 ( .A(n209), .B(n214), .Z(n207) );
  CIVX4 U1468 ( .A(n79), .Z(n1739) );
  CND2X1 U1469 ( .A(n666), .B(n683), .Z(n281) );
  CND2X1 U1470 ( .A(n631), .B(n633), .Z(n1566) );
  CND2X1 U1471 ( .A(n631), .B(n614), .Z(n1567) );
  CND2X1 U1472 ( .A(n633), .B(n614), .Z(n1568) );
  CND3X2 U1473 ( .A(n1566), .B(n1567), .C(n1568), .Z(n607) );
  CNR2XL U1474 ( .A(n36), .B(n1311), .Z(n1569) );
  CNR2XL U1475 ( .A(n1310), .B(n1621), .Z(n1570) );
  COR2X1 U1476 ( .A(n1569), .B(n1570), .Z(n1027) );
  COR2X2 U1477 ( .A(n77), .B(n1203), .Z(n1571) );
  CND2X2 U1478 ( .A(n1571), .B(n1572), .Z(n924) );
  CIVXL U1479 ( .A(a[8]), .Z(n1573) );
  CND2X1 U1480 ( .A(n1576), .B(n1577), .Z(n1579) );
  CIVXL U1481 ( .A(n1692), .Z(n1576) );
  CIVXL U1482 ( .A(n1738), .Z(n1577) );
  CIVX1 U1483 ( .A(n1739), .Z(n1738) );
  CND2X1 U1484 ( .A(a[14]), .B(n1726), .Z(n1582) );
  CIVX2 U1485 ( .A(a[14]), .Z(n1580) );
  CIVX2 U1486 ( .A(n1726), .Z(n1581) );
  CND2X1 U1487 ( .A(a[12]), .B(n1585), .Z(n1586) );
  CND2XL U1488 ( .A(n1584), .B(n1724), .Z(n1587) );
  CND2X1 U1489 ( .A(n1586), .B(n1587), .Z(n1447) );
  CIVX2 U1490 ( .A(a[12]), .Z(n1584) );
  CIVXL U1491 ( .A(n1724), .Z(n1585) );
  CND2X4 U1492 ( .A(n1447), .B(n58), .Z(n61) );
  CENXL U1493 ( .A(n1707), .B(n155), .Z(n1333) );
  CIVX2 U1494 ( .A(n12), .Z(n1705) );
  CENXL U1495 ( .A(n1724), .B(n152), .Z(n1232) );
  CENX4 U1496 ( .A(n1724), .B(a[14]), .Z(n66) );
  CNR2IX1 U1497 ( .B(n1691), .A(n105), .Z(n872) );
  CENX2 U1498 ( .A(n1689), .B(a[26]), .Z(n105) );
  CIVX2 U1499 ( .A(n1598), .Z(n1588) );
  CIVXL U1500 ( .A(n1588), .Z(n1589) );
  CIVXL U1501 ( .A(n1588), .Z(n1590) );
  CNIVX8 U1502 ( .A(n87), .Z(n1687) );
  CND2X4 U1503 ( .A(n1448), .B(n1624), .Z(n53) );
  CND2X1 U1504 ( .A(n1702), .B(a[4]), .Z(n1602) );
  COND2X1 U1505 ( .A(n18), .B(n1363), .C(n1362), .D(n15), .Z(n1077) );
  CENXL U1506 ( .A(n1695), .B(n109), .Z(n1135) );
  CIVXL U1507 ( .A(n109), .Z(n1464) );
  CENXL U1508 ( .A(n1690), .B(n109), .Z(n1138) );
  CENXL U1509 ( .A(n1693), .B(n109), .Z(n1137) );
  CENXL U1510 ( .A(n1676), .B(n109), .Z(n1136) );
  CND2IXL U1511 ( .B(n1691), .A(n109), .Z(n1139) );
  CENXL U1512 ( .A(n109), .B(a[30]), .Z(n114) );
  CENXL U1513 ( .A(n1721), .B(n155), .Z(n1252) );
  CENXL U1514 ( .A(n1721), .B(n154), .Z(n1253) );
  CENXL U1515 ( .A(n1721), .B(n1681), .Z(n1265) );
  CENXL U1516 ( .A(n1721), .B(n1679), .Z(n1267) );
  CENXL U1517 ( .A(n1721), .B(n152), .Z(n1255) );
  CENXL U1518 ( .A(n1721), .B(n1683), .Z(n1263) );
  CENXL U1519 ( .A(n1721), .B(n1676), .Z(n1271) );
  CENXL U1520 ( .A(n1721), .B(n142), .Z(n1261) );
  CENXL U1521 ( .A(n1721), .B(n146), .Z(n1259) );
  CENXL U1522 ( .A(n1721), .B(n150), .Z(n1257) );
  CENXL U1523 ( .A(n1721), .B(n1677), .Z(n1269) );
  COND2XL U1524 ( .A(n1156), .B(n95), .C(n1157), .D(n97), .Z(n881) );
  COND2XL U1525 ( .A(n1158), .B(n97), .C(n1157), .D(n95), .Z(n882) );
  COND2XL U1526 ( .A(n1158), .B(n95), .C(n1159), .D(n97), .Z(n883) );
  COND2XL U1527 ( .A(n1160), .B(n95), .C(n1161), .D(n97), .Z(n885) );
  COND2XL U1528 ( .A(n1561), .B(n1388), .C(n1696), .D(n1387), .Z(n1101) );
  COND2XL U1529 ( .A(n1561), .B(n1389), .C(n1696), .D(n1388), .Z(n1102) );
  COND2XL U1530 ( .A(n1561), .B(n1390), .C(n1696), .D(n1389), .Z(n1103) );
  COND2XL U1531 ( .A(n1675), .B(n1391), .C(n1696), .D(n1390), .Z(n1104) );
  COND2XL U1532 ( .A(n1561), .B(n1410), .C(n1696), .D(n1409), .Z(n1123) );
  COND2XL U1533 ( .A(n1561), .B(n1409), .C(n1696), .D(n1408), .Z(n1122) );
  COND2XL U1534 ( .A(n1675), .B(n1393), .C(n1696), .D(n1392), .Z(n1106) );
  COND2XL U1535 ( .A(n1675), .B(n1395), .C(n1696), .D(n1394), .Z(n1108) );
  COND2XL U1536 ( .A(n1675), .B(n1392), .C(n1696), .D(n1391), .Z(n1105) );
  COND2X1 U1537 ( .A(n1175), .B(n91), .C(n1174), .D(n1661), .Z(n898) );
  CND2X2 U1538 ( .A(n1443), .B(n89), .Z(n91) );
  CNIVX2 U1539 ( .A(n99), .Z(n1689) );
  CIVX1 U1540 ( .A(n55), .Z(n1725) );
  CIVX4 U1541 ( .A(n1725), .Z(n1724) );
  COND1X1 U1542 ( .A(n253), .B(n236), .C(n237), .Z(n235) );
  CND2IX2 U1543 ( .B(n1625), .A(n100), .Z(n102) );
  CENXL U1544 ( .A(n1680), .B(n1689), .Z(n1147) );
  CENXL U1545 ( .A(n1679), .B(n1689), .Z(n1148) );
  CENXL U1546 ( .A(n1678), .B(n1689), .Z(n1149) );
  CIVXL U1547 ( .A(n1689), .Z(n1466) );
  CND2IXL U1548 ( .B(n1691), .A(n1689), .Z(n1155) );
  COND1X1 U1549 ( .A(n217), .B(n209), .C(n210), .Z(n208) );
  CNR2X2 U1550 ( .A(n454), .B(n481), .Z(n209) );
  CND2XL U1551 ( .A(n879), .B(n1558), .Z(n1593) );
  CND2XL U1552 ( .A(n879), .B(n1077), .Z(n1594) );
  CND2XL U1553 ( .A(n1558), .B(n1077), .Z(n1595) );
  CND3X1 U1554 ( .A(n1593), .B(n1594), .C(n1595), .Z(n577) );
  CNR2XL U1555 ( .A(n1153), .B(n100), .Z(n1596) );
  CNR2XL U1556 ( .A(n102), .B(n1154), .Z(n1597) );
  COR2X1 U1557 ( .A(n1596), .B(n1597), .Z(n879) );
  CENXL U1558 ( .A(n1692), .B(n1689), .Z(n1153) );
  CENX4 U1559 ( .A(n1688), .B(a[24]), .Z(n100) );
  CENXL U1560 ( .A(n1690), .B(n1689), .Z(n1154) );
  CIVX2 U1561 ( .A(n30), .Z(n1714) );
  CANR1X1 U1562 ( .A(n220), .B(n207), .C(n208), .Z(n206) );
  COND1X1 U1563 ( .A(n231), .B(n225), .C(n226), .Z(n220) );
  CNR2X2 U1564 ( .A(n666), .B(n683), .Z(n280) );
  COND2XL U1565 ( .A(n27), .B(n1353), .C(n1352), .D(n1623), .Z(n1068) );
  CNIVX2 U1566 ( .A(n132), .Z(n1680) );
  CND2X1 U1567 ( .A(n1600), .B(n1601), .Z(n1603) );
  COND2XL U1568 ( .A(n27), .B(n1340), .C(n1339), .D(n1623), .Z(n1055) );
  COND2XL U1569 ( .A(n27), .B(n1332), .C(n1331), .D(n1623), .Z(n1047) );
  COND2XL U1570 ( .A(n27), .B(n1331), .C(n1330), .D(n1623), .Z(n1046) );
  COND2XL U1571 ( .A(n27), .B(n1345), .C(n1344), .D(n1623), .Z(n1060) );
  COND2XL U1572 ( .A(n27), .B(n1330), .C(n1329), .D(n1623), .Z(n1045) );
  COND2XL U1573 ( .A(n27), .B(n1352), .C(n1623), .D(n1351), .Z(n1067) );
  COND2XL U1574 ( .A(n27), .B(n1354), .C(n1623), .D(n1353), .Z(n1069) );
  CIVDX1 U1575 ( .A(n3), .Z0(n1599), .Z1(n1598) );
  CIVXL U1576 ( .A(n1702), .Z(n1600) );
  CANR1X1 U1577 ( .A(n1633), .B(n204), .C(n201), .Z(n199) );
  COND2X1 U1578 ( .A(n27), .B(n1336), .C(n1335), .D(n1623), .Z(n1051) );
  COND2XL U1579 ( .A(n77), .B(n1199), .C(n1198), .D(n1557), .Z(n920) );
  COND2XL U1580 ( .A(n77), .B(n1200), .C(n1557), .D(n1199), .Z(n921) );
  COND2XL U1581 ( .A(n44), .B(n1293), .C(n1292), .D(n42), .Z(n1010) );
  COND2X1 U1582 ( .A(n27), .B(n1333), .C(n1332), .D(n1623), .Z(n1048) );
  COND2XL U1583 ( .A(n77), .B(n1198), .C(n1557), .D(n1197), .Z(n919) );
  COND2X1 U1584 ( .A(n27), .B(n1351), .C(n1350), .D(n1623), .Z(n1066) );
  COND2XL U1585 ( .A(n27), .B(n1347), .C(n1346), .D(n1623), .Z(n1062) );
  COND2XL U1586 ( .A(n36), .B(n1325), .C(n1621), .D(n1324), .Z(n1041) );
  CND2IXL U1587 ( .B(n1691), .A(n1706), .Z(n1355) );
  CNR2IX1 U1588 ( .B(n1691), .A(n1623), .Z(n1070) );
  COND2XL U1589 ( .A(n27), .B(n1334), .C(n1333), .D(n1623), .Z(n1049) );
  CNIVX4 U1590 ( .A(n126), .Z(n1677) );
  CND2X4 U1591 ( .A(n1602), .B(n1603), .Z(n1623) );
  CIVXL U1592 ( .A(a[4]), .Z(n1601) );
  COND2X1 U1593 ( .A(n27), .B(n1341), .C(n1340), .D(n1623), .Z(n1056) );
  CND2IX4 U1594 ( .B(n1622), .A(n1623), .Z(n27) );
  COND2XL U1595 ( .A(n27), .B(n1553), .C(n1355), .D(n1623), .Z(n858) );
  COND2X1 U1596 ( .A(n53), .B(n1267), .C(n1624), .D(n1266), .Z(n985) );
  COND2X1 U1597 ( .A(n1190), .B(n1657), .C(n1191), .D(n85), .Z(n913) );
  COND2X1 U1598 ( .A(n1188), .B(n1657), .C(n1189), .D(n85), .Z(n911) );
  CIVX4 U1599 ( .A(n71), .Z(n1734) );
  CANR1X1 U1600 ( .A(n212), .B(n232), .C(n213), .Z(n211) );
  CNR2IX1 U1601 ( .B(n1691), .A(n110), .Z(n866) );
  COND2XL U1602 ( .A(n36), .B(n1309), .C(n1308), .D(n1621), .Z(n1025) );
  COND2XL U1603 ( .A(n36), .B(n1319), .C(n1621), .D(n1318), .Z(n1035) );
  CND2X1 U1604 ( .A(n1609), .B(n1610), .Z(n1612) );
  CIVX1 U1605 ( .A(n233), .Z(n232) );
  CIVXL U1606 ( .A(n209), .Z(n381) );
  CND2XL U1607 ( .A(n1729), .B(a[18]), .Z(n1606) );
  CND2X1 U1608 ( .A(n1604), .B(n1605), .Z(n1607) );
  CND2X2 U1609 ( .A(n1606), .B(n1607), .Z(n1657) );
  CIVXL U1610 ( .A(n1729), .Z(n1604) );
  CIVXL U1611 ( .A(a[18]), .Z(n1605) );
  CANR1X1 U1612 ( .A(n304), .B(n1636), .C(n297), .Z(n295) );
  CIVX2 U1613 ( .A(n1553), .Z(n1707) );
  CND2IXL U1614 ( .B(n1691), .A(n55), .Z(n1251) );
  COND2X1 U1615 ( .A(n36), .B(n1322), .C(n1321), .D(n1621), .Z(n1038) );
  CNR2IXL U1616 ( .B(n1691), .A(n1621), .Z(n1042) );
  CIVXL U1617 ( .A(n21), .Z(n1609) );
  COAN1XL U1618 ( .A(n288), .B(n271), .C(n272), .Z(n1608) );
  CND2X4 U1619 ( .A(n1611), .B(n1612), .Z(n1621) );
  CIVXL U1620 ( .A(a[6]), .Z(n1610) );
  COND2XL U1621 ( .A(n36), .B(n1301), .C(n1300), .D(n1621), .Z(n1017) );
  CND2X4 U1622 ( .A(n1450), .B(n1621), .Z(n36) );
  CAN2X1 U1623 ( .A(n1633), .B(n203), .Z(n1617) );
  CND2X1 U1624 ( .A(n482), .B(n507), .Z(n217) );
  CIVX1 U1625 ( .A(n264), .Z(n266) );
  CIVX1 U1626 ( .A(n259), .Z(n1627) );
  CND2XL U1627 ( .A(n392), .B(n292), .Z(n179) );
  CANR1XL U1628 ( .A(n376), .B(n1646), .C(n373), .Z(n371) );
  CANR1XL U1629 ( .A(n368), .B(n1647), .C(n365), .Z(n363) );
  CENX1 U1630 ( .A(n193), .B(n368), .Z(product[4]) );
  CND2XL U1631 ( .A(n407), .B(n370), .Z(n194) );
  CND2X1 U1632 ( .A(n1050), .B(n958), .Z(n1668) );
  COND2XL U1633 ( .A(n27), .B(n1338), .C(n1337), .D(n1623), .Z(n1053) );
  COND2X1 U1634 ( .A(n85), .B(n1184), .C(n1183), .D(n1657), .Z(n906) );
  COND2XL U1635 ( .A(n1675), .B(n1415), .C(n1696), .D(n1414), .Z(n1128) );
  CND2X1 U1636 ( .A(n1614), .B(a[16]), .Z(n1630) );
  CIVX2 U1637 ( .A(a[16]), .Z(n1629) );
  CNIVX1 U1638 ( .A(n120), .Z(n1692) );
  CNIVX1 U1639 ( .A(n144), .Z(n1685) );
  COND1XL U1640 ( .A(n205), .B(n1592), .C(n1560), .Z(n1613) );
  CNIVX4 U1641 ( .A(n63), .Z(n1614) );
  CENXL U1642 ( .A(n1615), .B(n227), .Z(product[27]) );
  CAN2XL U1643 ( .A(n383), .B(n226), .Z(n1615) );
  CENXL U1644 ( .A(n1616), .B(n218), .Z(product[28]) );
  CEOXL U1645 ( .A(n168), .B(n211), .Z(product[29]) );
  CEOXL U1646 ( .A(n1613), .B(n1617), .Z(product[30]) );
  COND1X1 U1647 ( .A(n309), .B(n321), .C(n310), .Z(n308) );
  CANR1X1 U1648 ( .A(n308), .B(n289), .C(n290), .Z(n288) );
  CNR2X2 U1649 ( .A(n508), .B(n533), .Z(n225) );
  CIVX1 U1650 ( .A(n299), .Z(n297) );
  CND2XL U1651 ( .A(n1636), .B(n394), .Z(n294) );
  CND2XL U1652 ( .A(n1635), .B(n276), .Z(n176) );
  CEOXL U1653 ( .A(n176), .B(n277), .Z(product[21]) );
  CEOXL U1654 ( .A(n177), .B(n282), .Z(product[20]) );
  CEOXL U1655 ( .A(n182), .B(n315), .Z(product[15]) );
  CND2XL U1656 ( .A(n1638), .B(n314), .Z(n182) );
  CEOXL U1657 ( .A(n181), .B(n307), .Z(product[16]) );
  CND2XL U1658 ( .A(n394), .B(n302), .Z(n181) );
  COND1XL U1659 ( .A(n252), .B(n1608), .C(n253), .Z(n251) );
  CND2XL U1660 ( .A(n254), .B(n1639), .Z(n243) );
  CND2XL U1661 ( .A(n391), .B(n286), .Z(n178) );
  CND2XL U1662 ( .A(n1637), .B(n319), .Z(n183) );
  CANR1X1 U1663 ( .A(n330), .B(n322), .C(n323), .Z(n321) );
  CNR2XL U1664 ( .A(n324), .B(n327), .Z(n322) );
  CANR1X1 U1665 ( .A(n352), .B(n344), .C(n345), .Z(n343) );
  COND1X1 U1666 ( .A(n331), .B(n343), .C(n332), .Z(n330) );
  CND2XL U1667 ( .A(n1641), .B(n1642), .Z(n331) );
  CND2XL U1668 ( .A(n702), .B(n717), .Z(n292) );
  CND2XL U1669 ( .A(n402), .B(n350), .Z(n189) );
  CND2XL U1670 ( .A(n1641), .B(n336), .Z(n186) );
  CND2XL U1671 ( .A(n398), .B(n328), .Z(n185) );
  CEOXL U1672 ( .A(n185), .B(n329), .Z(product[12]) );
  CND2XL U1673 ( .A(n1642), .B(n341), .Z(n187) );
  CANR1X1 U1674 ( .A(n360), .B(n1648), .C(n357), .Z(n355) );
  CENXL U1675 ( .A(n1665), .B(n199), .Z(product[31]) );
  CND2XL U1676 ( .A(n425), .B(n410), .Z(n198) );
  CND2XL U1677 ( .A(n814), .B(n821), .Z(n347) );
  CND2XL U1678 ( .A(n403), .B(n354), .Z(n190) );
  CEOXL U1679 ( .A(n190), .B(n355), .Z(product[7]) );
  CENXL U1680 ( .A(n191), .B(n360), .Z(product[6]) );
  CND2XL U1681 ( .A(n1648), .B(n359), .Z(n191) );
  CND2XL U1682 ( .A(n774), .B(n785), .Z(n325) );
  CND2XL U1683 ( .A(n1646), .B(n375), .Z(n195) );
  CND2XL U1684 ( .A(n1647), .B(n367), .Z(n193) );
  CEOXL U1685 ( .A(n371), .B(n194), .Z(product[3]) );
  CND2XL U1686 ( .A(n405), .B(n362), .Z(n192) );
  CEOXL U1687 ( .A(n363), .B(n192), .Z(product[5]) );
  CND3X1 U1688 ( .A(n1662), .B(n1663), .C(n1664), .Z(n573) );
  CND3X1 U1689 ( .A(n1666), .B(n1667), .C(n1668), .Z(n595) );
  CND2XL U1690 ( .A(n844), .B(n1129), .Z(n370) );
  COR2XL U1691 ( .A(n1131), .B(n860), .Z(n1618) );
  CNR2IXL U1692 ( .B(n1691), .A(n1557), .Z(n932) );
  COND2XL U1693 ( .A(n77), .B(n1206), .C(n1557), .D(n1205), .Z(n927) );
  COND2XL U1694 ( .A(n77), .B(n1201), .C(n1200), .D(n1557), .Z(n922) );
  CNIVXL U1695 ( .A(n124), .Z(n1695) );
  CEO3X1 U1696 ( .A(n449), .B(n443), .C(n445), .Z(n417) );
  CEO3X1 U1697 ( .A(n423), .B(n421), .C(n420), .Z(n416) );
  CEO3XL U1698 ( .A(n867), .B(n917), .C(n971), .Z(n420) );
  CEO3XL U1699 ( .A(n881), .B(n933), .C(n993), .Z(n423) );
  CENX1 U1700 ( .A(a[18]), .B(n1736), .Z(n1619) );
  CND2IX4 U1701 ( .B(n1620), .A(n15), .Z(n18) );
  CENX1 U1702 ( .A(a[2]), .B(n1702), .Z(n1620) );
  CENX4 U1703 ( .A(n1721), .B(a[12]), .Z(n58) );
  CENX4 U1704 ( .A(n1716), .B(a[10]), .Z(n1624) );
  CNIVX4 U1705 ( .A(n130), .Z(n1679) );
  CND2XL U1706 ( .A(n1438), .B(n114), .Z(n115) );
  CNIVX3 U1707 ( .A(n128), .Z(n1678) );
  CND2X1 U1708 ( .A(n266), .B(n1632), .Z(n1626) );
  CIVXL U1709 ( .A(n253), .Z(n255) );
  CNR2IXL U1710 ( .B(n219), .A(n214), .Z(n212) );
  COND1XL U1711 ( .A(n205), .B(n1592), .C(n206), .Z(n204) );
  CND2XL U1712 ( .A(n381), .B(n210), .Z(n168) );
  CND2X1 U1713 ( .A(n1632), .B(n388), .Z(n252) );
  CND2XL U1714 ( .A(n278), .B(n1635), .Z(n271) );
  CENX1 U1715 ( .A(n232), .B(n171), .Z(product[26]) );
  CANR1X1 U1716 ( .A(n270), .B(n234), .C(n235), .Z(n233) );
  CANR1XL U1717 ( .A(n1639), .B(n255), .C(n248), .Z(n244) );
  CENX1 U1718 ( .A(n262), .B(n174), .Z(product[23]) );
  COND1XL U1719 ( .A(n263), .B(n1608), .C(n264), .Z(n262) );
  CENX1 U1720 ( .A(n320), .B(n183), .Z(product[14]) );
  CENX1 U1721 ( .A(n300), .B(n180), .Z(product[17]) );
  CND2X1 U1722 ( .A(n1636), .B(n299), .Z(n180) );
  COND1XL U1723 ( .A(n301), .B(n307), .C(n302), .Z(n300) );
  CENX1 U1724 ( .A(n287), .B(n178), .Z(product[19]) );
  COND1XL U1725 ( .A(n243), .B(n1608), .C(n244), .Z(n242) );
  CND2X1 U1726 ( .A(n390), .B(n281), .Z(n177) );
  CANR1XL U1727 ( .A(n391), .B(n287), .C(n284), .Z(n282) );
  CEOXL U1728 ( .A(n175), .B(n1608), .Z(product[22]) );
  CANR1XL U1729 ( .A(n1637), .B(n320), .C(n317), .Z(n315) );
  COR2X1 U1730 ( .A(n604), .B(n625), .Z(n1632) );
  CND2X1 U1731 ( .A(n604), .B(n625), .Z(n261) );
  CND2X1 U1732 ( .A(n426), .B(n453), .Z(n203) );
  COR2X1 U1733 ( .A(n426), .B(n453), .Z(n1633) );
  CENX1 U1734 ( .A(n606), .B(n1634), .Z(n604) );
  CENX1 U1735 ( .A(n608), .B(n627), .Z(n1634) );
  COND1XL U1736 ( .A(n328), .B(n324), .C(n325), .Z(n323) );
  CNR2X1 U1737 ( .A(n346), .B(n349), .Z(n344) );
  COND1XL U1738 ( .A(n350), .B(n346), .C(n347), .Z(n345) );
  CANR1XL U1739 ( .A(n339), .B(n1641), .C(n334), .Z(n332) );
  CENX1 U1740 ( .A(n188), .B(n348), .Z(product[9]) );
  CND2X1 U1741 ( .A(n401), .B(n347), .Z(n188) );
  COND1XL U1742 ( .A(n349), .B(n351), .C(n350), .Z(n348) );
  CENX1 U1743 ( .A(n342), .B(n187), .Z(product[10]) );
  CENX1 U1744 ( .A(n326), .B(n184), .Z(product[13]) );
  CND2X1 U1745 ( .A(n397), .B(n325), .Z(n184) );
  COND1XL U1746 ( .A(n327), .B(n329), .C(n328), .Z(n326) );
  CNR2X1 U1747 ( .A(n684), .B(n701), .Z(n285) );
  CNR2X1 U1748 ( .A(n734), .B(n747), .Z(n301) );
  COR2X1 U1749 ( .A(n646), .B(n665), .Z(n1635) );
  CEOX1 U1750 ( .A(n351), .B(n189), .Z(product[8]) );
  CEOX1 U1751 ( .A(n186), .B(n337), .Z(product[11]) );
  CANR1XL U1752 ( .A(n1642), .B(n342), .C(n339), .Z(n337) );
  COR2X1 U1753 ( .A(n718), .B(n733), .Z(n1636) );
  CND2X1 U1754 ( .A(n684), .B(n701), .Z(n286) );
  CNR2X1 U1755 ( .A(n534), .B(n557), .Z(n230) );
  COR2X1 U1756 ( .A(n762), .B(n773), .Z(n1637) );
  CND2X1 U1757 ( .A(n734), .B(n747), .Z(n302) );
  COR2X1 U1758 ( .A(n582), .B(n603), .Z(n1639) );
  CND2X1 U1759 ( .A(n762), .B(n773), .Z(n319) );
  CND2X1 U1760 ( .A(n748), .B(n761), .Z(n314) );
  CND2X1 U1761 ( .A(n646), .B(n665), .Z(n276) );
  CND2X1 U1762 ( .A(n718), .B(n733), .Z(n299) );
  CND2X1 U1763 ( .A(n626), .B(n645), .Z(n264) );
  COR2X1 U1764 ( .A(n581), .B(n558), .Z(n1640) );
  CND2X1 U1765 ( .A(n558), .B(n581), .Z(n241) );
  COND1XL U1766 ( .A(n371), .B(n369), .C(n370), .Z(n368) );
  COND1XL U1767 ( .A(n363), .B(n361), .C(n362), .Z(n360) );
  COND1XL U1768 ( .A(n353), .B(n355), .C(n354), .Z(n352) );
  CAN2X1 U1769 ( .A(n1643), .B(n198), .Z(n1665) );
  CNR2X1 U1770 ( .A(n822), .B(n827), .Z(n349) );
  CNR2X1 U1771 ( .A(n786), .B(n795), .Z(n327) );
  CNR2X1 U1772 ( .A(n774), .B(n785), .Z(n324) );
  CNR2X1 U1773 ( .A(n814), .B(n821), .Z(n346) );
  COR2X1 U1774 ( .A(n796), .B(n805), .Z(n1641) );
  COR2X1 U1775 ( .A(n806), .B(n813), .Z(n1642) );
  CND2X1 U1776 ( .A(n822), .B(n827), .Z(n350) );
  CND2X1 U1777 ( .A(n786), .B(n795), .Z(n328) );
  CND2X1 U1778 ( .A(n806), .B(n813), .Z(n341) );
  CND2X1 U1779 ( .A(n796), .B(n805), .Z(n336) );
  COR2X1 U1780 ( .A(n425), .B(n410), .Z(n1643) );
  CENX1 U1781 ( .A(n195), .B(n376), .Z(product[2]) );
  CENX1 U1782 ( .A(n1694), .B(n1712), .Z(n1322) );
  CENX1 U1783 ( .A(n1694), .B(n1590), .Z(n1415) );
  CENX1 U1784 ( .A(n1694), .B(n1704), .Z(n1382) );
  CENX1 U1785 ( .A(n1694), .B(n1717), .Z(n1295) );
  CENX1 U1786 ( .A(n1694), .B(n1722), .Z(n1270) );
  CENX1 U1787 ( .A(n1694), .B(n1737), .Z(n1190) );
  CENX1 U1788 ( .A(n1694), .B(n1554), .Z(n1351) );
  CENX1 U1789 ( .A(n1694), .B(n1731), .Z(n1207) );
  CNR2X1 U1790 ( .A(n828), .B(n833), .Z(n353) );
  CNR2X1 U1791 ( .A(n844), .B(n1129), .Z(n369) );
  CNR2X1 U1792 ( .A(n838), .B(n841), .Z(n361) );
  CND3XL U1793 ( .A(n1669), .B(n1670), .C(n1671), .Z(n589) );
  CENX1 U1794 ( .A(n1644), .B(n596), .Z(n590) );
  CENX1 U1795 ( .A(n1645), .B(n1049), .Z(n574) );
  CENX1 U1796 ( .A(n977), .B(n939), .Z(n1645) );
  CND2X1 U1797 ( .A(n1131), .B(n860), .Z(n378) );
  CND2X1 U1798 ( .A(n1130), .B(n1100), .Z(n375) );
  CND2X1 U1799 ( .A(n842), .B(n843), .Z(n367) );
  CND2X1 U1800 ( .A(n834), .B(n837), .Z(n359) );
  CND2X1 U1801 ( .A(n838), .B(n841), .Z(n362) );
  CND2X1 U1802 ( .A(n828), .B(n833), .Z(n354) );
  COR2X1 U1803 ( .A(n1130), .B(n1100), .Z(n1646) );
  COR2X1 U1804 ( .A(n842), .B(n843), .Z(n1647) );
  COR2X1 U1805 ( .A(n834), .B(n837), .Z(n1648) );
  CIVX2 U1806 ( .A(n1599), .Z(n1698) );
  CENX1 U1807 ( .A(n151), .B(n1726), .Z(n1212) );
  CENX1 U1808 ( .A(n1735), .B(n1676), .Z(n1191) );
  CENX1 U1809 ( .A(n1702), .B(n1676), .Z(n1383) );
  CENX1 U1810 ( .A(n1710), .B(n1676), .Z(n1323) );
  CENX1 U1811 ( .A(n1685), .B(n1711), .Z(n1312) );
  CENX1 U1812 ( .A(n1614), .B(n1679), .Z(n1223) );
  CENX1 U1813 ( .A(n1702), .B(n1683), .Z(n1375) );
  CENX1 U1814 ( .A(n1711), .B(n1681), .Z(n1317) );
  CENX1 U1815 ( .A(n1709), .B(n151), .Z(n1308) );
  CENX1 U1816 ( .A(n1735), .B(n1679), .Z(n1187) );
  CENX1 U1817 ( .A(n1709), .B(n153), .Z(n1306) );
  CENX1 U1818 ( .A(n151), .B(n1717), .Z(n1281) );
  CENX1 U1819 ( .A(n1554), .B(n151), .Z(n1337) );
  CENX1 U1820 ( .A(n1701), .B(n1679), .Z(n1379) );
  CENX1 U1821 ( .A(n1700), .B(n1681), .Z(n1377) );
  CENX1 U1822 ( .A(n153), .B(n1722), .Z(n1254) );
  CENX1 U1823 ( .A(n1701), .B(n1677), .Z(n1381) );
  CENX1 U1824 ( .A(n1690), .B(n1589), .Z(n1418) );
  CENX1 U1825 ( .A(n1682), .B(n1704), .Z(n1376) );
  CENX1 U1826 ( .A(n1678), .B(n1709), .Z(n1320) );
  CENX1 U1827 ( .A(n1680), .B(n1711), .Z(n1318) );
  CENX1 U1828 ( .A(n1589), .B(n151), .Z(n1401) );
  CENX1 U1829 ( .A(n151), .B(n1722), .Z(n1256) );
  CENX1 U1830 ( .A(n1682), .B(n1738), .Z(n1184) );
  CENX1 U1831 ( .A(n1680), .B(n1737), .Z(n1186) );
  CENX1 U1832 ( .A(n1697), .B(n1679), .Z(n1412) );
  CENX1 U1833 ( .A(n1680), .B(n1704), .Z(n1378) );
  CENX1 U1834 ( .A(n1678), .B(n1704), .Z(n1380) );
  CENX1 U1835 ( .A(n1678), .B(n1737), .Z(n1188) );
  CENX1 U1836 ( .A(n1694), .B(n1688), .Z(n1162) );
  CENX1 U1837 ( .A(n1700), .B(n151), .Z(n1368) );
  CENX1 U1838 ( .A(n1726), .B(n1676), .Z(n1227) );
  CENX1 U1839 ( .A(n1727), .B(n1683), .Z(n1219) );
  CENX1 U1840 ( .A(n1684), .B(n1717), .Z(n1287) );
  CENX1 U1841 ( .A(n1684), .B(n1738), .Z(n1182) );
  CENX1 U1842 ( .A(n1685), .B(n1737), .Z(n1180) );
  CIVX2 U1843 ( .A(n1723), .Z(n1722) );
  CENX1 U1844 ( .A(n1690), .B(n1738), .Z(n1193) );
  CENX1 U1845 ( .A(n1699), .B(n153), .Z(n1366) );
  CENX1 U1846 ( .A(n1715), .B(n153), .Z(n1279) );
  CENX1 U1847 ( .A(n1678), .B(n1731), .Z(n1205) );
  CENX1 U1848 ( .A(n1680), .B(n1732), .Z(n1203) );
  CIVX2 U1849 ( .A(n1599), .Z(n1697) );
  CENX1 U1850 ( .A(n1682), .B(n1688), .Z(n1156) );
  CENX1 U1851 ( .A(n1686), .B(n1722), .Z(n1258) );
  CNR2IXL U1852 ( .B(n1691), .A(n15), .Z(n1100) );
  CENX1 U1853 ( .A(n1736), .B(n1677), .Z(n1189) );
  CENX1 U1854 ( .A(n1676), .B(n1688), .Z(n1163) );
  CENX1 U1855 ( .A(n1679), .B(n1688), .Z(n1159) );
  CENX1 U1856 ( .A(n1677), .B(n1688), .Z(n1161) );
  CENX1 U1857 ( .A(n1681), .B(n1688), .Z(n1157) );
  CENX1 U1858 ( .A(n1710), .B(n1677), .Z(n1321) );
  CENX1 U1859 ( .A(n1706), .B(n1677), .Z(n1350) );
  CENX1 U1860 ( .A(n1710), .B(n1679), .Z(n1319) );
  CENX1 U1861 ( .A(n1554), .B(n1679), .Z(n1348) );
  CENX1 U1862 ( .A(n1711), .B(n1686), .Z(n1310) );
  CENX1 U1863 ( .A(n1711), .B(n1683), .Z(n1315) );
  CENX1 U1864 ( .A(n1715), .B(n1681), .Z(n1290) );
  CENX1 U1865 ( .A(n1708), .B(n1683), .Z(n1344) );
  CENX1 U1866 ( .A(n1686), .B(n1717), .Z(n1283) );
  CENX1 U1867 ( .A(n1736), .B(n1683), .Z(n1183) );
  CENX1 U1868 ( .A(n1736), .B(n1681), .Z(n1185) );
  CENX1 U1869 ( .A(n1715), .B(n1676), .Z(n1296) );
  CENX1 U1870 ( .A(n1717), .B(n1677), .Z(n1294) );
  CENX1 U1871 ( .A(n1715), .B(n1679), .Z(n1292) );
  CENX1 U1872 ( .A(n1698), .B(n1676), .Z(n1416) );
  CENX1 U1873 ( .A(n1698), .B(n1677), .Z(n1414) );
  CENX1 U1874 ( .A(n1698), .B(n1683), .Z(n1408) );
  CENX1 U1875 ( .A(n1698), .B(n1684), .Z(n1407) );
  CENX1 U1876 ( .A(n1682), .B(n1722), .Z(n1264) );
  CENX1 U1877 ( .A(n1698), .B(n1685), .Z(n1405) );
  CENX1 U1878 ( .A(n1685), .B(n1717), .Z(n1285) );
  CENX1 U1879 ( .A(n1682), .B(n1717), .Z(n1289) );
  CENX1 U1880 ( .A(n1678), .B(n1722), .Z(n1268) );
  CENX1 U1881 ( .A(n1698), .B(n1686), .Z(n1403) );
  CENX1 U1882 ( .A(n1685), .B(n1722), .Z(n1260) );
  CENX1 U1883 ( .A(n1680), .B(n1717), .Z(n1291) );
  CENX1 U1884 ( .A(n1682), .B(n1712), .Z(n1316) );
  CENX1 U1885 ( .A(n1678), .B(n1717), .Z(n1293) );
  CENX1 U1886 ( .A(n1678), .B(n1589), .Z(n1413) );
  CENX1 U1887 ( .A(n1698), .B(n1681), .Z(n1410) );
  CENX1 U1888 ( .A(n1680), .B(n1590), .Z(n1411) );
  CENX1 U1889 ( .A(n1678), .B(n1554), .Z(n1349) );
  CENX1 U1890 ( .A(n1682), .B(n1590), .Z(n1409) );
  CENX1 U1891 ( .A(n1684), .B(n1722), .Z(n1262) );
  CENX1 U1892 ( .A(n1680), .B(n1722), .Z(n1266) );
  CENX1 U1893 ( .A(n1678), .B(n1688), .Z(n1160) );
  CENX1 U1894 ( .A(n1680), .B(n1688), .Z(n1158) );
  CENX1 U1895 ( .A(n1706), .B(n1676), .Z(n1352) );
  CENX1 U1896 ( .A(n1708), .B(n1685), .Z(n1341) );
  CENX1 U1897 ( .A(n1715), .B(n1683), .Z(n1288) );
  CENX1 U1898 ( .A(n1554), .B(n1681), .Z(n1346) );
  CENX1 U1899 ( .A(n1682), .B(n1727), .Z(n1220) );
  CENX1 U1900 ( .A(n1684), .B(n1727), .Z(n1218) );
  CENX1 U1901 ( .A(n1691), .B(n1727), .Z(n1229) );
  CENX1 U1902 ( .A(n1690), .B(n1717), .Z(n1298) );
  CENX1 U1903 ( .A(n1690), .B(n1712), .Z(n1325) );
  CENX1 U1904 ( .A(n1690), .B(n1688), .Z(n1165) );
  CENX1 U1905 ( .A(n1687), .B(n1677), .Z(n1174) );
  CENX1 U1906 ( .A(n1729), .B(n1676), .Z(n1208) );
  CENX1 U1907 ( .A(n1729), .B(n1679), .Z(n1204) );
  CENX1 U1908 ( .A(n1730), .B(n1677), .Z(n1206) );
  CENX1 U1909 ( .A(n1730), .B(n1683), .Z(n1200) );
  CENX1 U1910 ( .A(n1730), .B(n1681), .Z(n1202) );
  CENX1 U1911 ( .A(n1678), .B(n1687), .Z(n1173) );
  CENX1 U1912 ( .A(n1685), .B(n1727), .Z(n1216) );
  CENX1 U1913 ( .A(n1686), .B(n1727), .Z(n1214) );
  CENX1 U1914 ( .A(n1684), .B(n1733), .Z(n1199) );
  CENX1 U1915 ( .A(n1682), .B(n1732), .Z(n1201) );
  CENX1 U1916 ( .A(n1685), .B(n1733), .Z(n1197) );
  CIVX2 U1917 ( .A(n1734), .Z(n1730) );
  CIVX2 U1918 ( .A(n1734), .Z(n1732) );
  CENX1 U1919 ( .A(n1690), .B(n1700), .Z(n1385) );
  CENX1 U1920 ( .A(n1691), .B(n1732), .Z(n1210) );
  CNIVX1 U1921 ( .A(n926), .Z(n1654) );
  CNR2IXL U1922 ( .B(n1691), .A(n58), .Z(n970) );
  CNR2IXL U1923 ( .B(n1691), .A(n95), .Z(n890) );
  CENX1 U1924 ( .A(n1690), .B(n1722), .Z(n1273) );
  CNR2IXL U1925 ( .B(n1691), .A(n42), .Z(n1016) );
  CNR2IXL U1926 ( .B(n1691), .A(n1624), .Z(n992) );
  CEOX1 U1927 ( .A(n845), .B(n873), .Z(n424) );
  CIVX2 U1928 ( .A(n1734), .Z(n1731) );
  CNR2IXL U1929 ( .B(n1691), .A(n1696), .Z(product[0]) );
  CENX1 U1930 ( .A(n1710), .B(n150), .Z(n1309) );
  CENX1 U1931 ( .A(n1703), .B(n150), .Z(n1369) );
  CENX1 U1932 ( .A(n1711), .B(n142), .Z(n1313) );
  CENX1 U1933 ( .A(n1703), .B(n146), .Z(n1371) );
  CENX1 U1934 ( .A(n1701), .B(n142), .Z(n1373) );
  CENX1 U1935 ( .A(n1700), .B(n156), .Z(n1363) );
  CENX1 U1936 ( .A(n1710), .B(n156), .Z(n1303) );
  CENX1 U1937 ( .A(n1700), .B(b[25]), .Z(n1360) );
  CENX1 U1938 ( .A(n1700), .B(n157), .Z(n1362) );
  CENX1 U1939 ( .A(n1699), .B(b[27]), .Z(n1358) );
  CENX1 U1940 ( .A(n1717), .B(n156), .Z(n1276) );
  CENX1 U1941 ( .A(n1699), .B(b[28]), .Z(n1357) );
  CENX1 U1942 ( .A(n1697), .B(n154), .Z(n1398) );
  CENX1 U1943 ( .A(n1697), .B(n157), .Z(n1395) );
  CENX1 U1944 ( .A(n1697), .B(b[28]), .Z(n1390) );
  CENX1 U1945 ( .A(n1697), .B(b[27]), .Z(n1391) );
  CENX1 U1946 ( .A(n1697), .B(b[25]), .Z(n1393) );
  CENX1 U1947 ( .A(n1697), .B(b[26]), .Z(n1392) );
  CENX1 U1948 ( .A(n1697), .B(b[30]), .Z(n1388) );
  CENX1 U1949 ( .A(n104), .B(a[28]), .Z(n110) );
  CNIVX1 U1950 ( .A(n148), .Z(n1686) );
  CENX1 U1951 ( .A(n1701), .B(n154), .Z(n1365) );
  CENX1 U1952 ( .A(n1554), .B(b[27]), .Z(n1327) );
  CENX1 U1953 ( .A(n1709), .B(b[25]), .Z(n1300) );
  CENX1 U1954 ( .A(n1715), .B(n157), .Z(n1275) );
  CENX1 U1955 ( .A(n1690), .B(n113), .Z(n1133) );
  CENX1 U1956 ( .A(n1693), .B(n113), .Z(n1132) );
  CENX1 U1957 ( .A(n1701), .B(n152), .Z(n1367) );
  CENX1 U1958 ( .A(n1614), .B(n146), .Z(n1215) );
  CENX1 U1959 ( .A(n1727), .B(n142), .Z(n1217) );
  CENX1 U1960 ( .A(n1614), .B(n150), .Z(n1213) );
  CENX1 U1961 ( .A(n1735), .B(n142), .Z(n1181) );
  CENX1 U1962 ( .A(n1678), .B(n104), .Z(n1140) );
  CENX1 U1963 ( .A(n1554), .B(n150), .Z(n1338) );
  CENX1 U1964 ( .A(n1709), .B(n157), .Z(n1302) );
  CENX1 U1965 ( .A(n1710), .B(n154), .Z(n1305) );
  CENX1 U1966 ( .A(n1706), .B(n142), .Z(n1342) );
  CENX1 U1967 ( .A(n1554), .B(n157), .Z(n1331) );
  CENX1 U1968 ( .A(n1709), .B(b[24]), .Z(n1301) );
  CENX1 U1969 ( .A(n1676), .B(n104), .Z(n1143) );
  CENX1 U1970 ( .A(n1677), .B(n104), .Z(n1141) );
  CENX1 U1971 ( .A(n1698), .B(n142), .Z(n1406) );
  CENX1 U1972 ( .A(n1698), .B(n150), .Z(n1402) );
  CENX1 U1973 ( .A(n1698), .B(n146), .Z(n1404) );
  CENX1 U1974 ( .A(n1695), .B(n104), .Z(n1142) );
  CENX1 U1975 ( .A(n1708), .B(b[24]), .Z(n1330) );
  CENX1 U1976 ( .A(n1715), .B(n154), .Z(n1278) );
  CENX1 U1977 ( .A(n1698), .B(b[31]), .Z(n1387) );
  CENX1 U1978 ( .A(n1730), .B(n142), .Z(n1198) );
  CENX1 U1979 ( .A(n1729), .B(n146), .Z(n1196) );
  CENX1 U1980 ( .A(n1554), .B(b[25]), .Z(n1329) );
  CENX1 U1981 ( .A(n1554), .B(b[26]), .Z(n1328) );
  CENX1 U1982 ( .A(n1714), .B(a[8]), .Z(n1656) );
  CNIVX4 U1983 ( .A(n122), .Z(n1676) );
  CND2X1 U1984 ( .A(n1439), .B(n110), .Z(n112) );
  CEOXL U1985 ( .A(a[28]), .B(n109), .Z(n1439) );
  CIVX2 U1986 ( .A(n39), .Z(n1719) );
  CNIVX2 U1987 ( .A(n134), .Z(n1681) );
  CNIVXL U1988 ( .A(n120), .Z(n1693) );
  CEOX1 U1989 ( .A(a[30]), .B(n113), .Z(n1438) );
  CIVX1 U1990 ( .A(n900), .Z(n1650) );
  CIVX2 U1991 ( .A(n1650), .Z(n1651) );
  CENX1 U1992 ( .A(n1697), .B(b[24]), .Z(n1394) );
  CENX1 U1993 ( .A(n1697), .B(n156), .Z(n1396) );
  CENX1 U1994 ( .A(n1697), .B(n153), .Z(n1399) );
  COND2XL U1995 ( .A(n69), .B(n1213), .C(n66), .D(n1212), .Z(n933) );
  COND2XL U1996 ( .A(n69), .B(n1215), .C(n66), .D(n1214), .Z(n935) );
  COND2XL U1997 ( .A(n69), .B(n1214), .C(n1213), .D(n66), .Z(n934) );
  COND2XL U1998 ( .A(n69), .B(n1217), .C(n66), .D(n1216), .Z(n937) );
  CNR2IXL U1999 ( .B(n1691), .A(n66), .Z(n950) );
  COND2XL U2000 ( .A(n69), .B(n1218), .C(n1217), .D(n66), .Z(n938) );
  COND2XL U2001 ( .A(n69), .B(n1229), .C(n66), .D(n1228), .Z(n949) );
  COND2XL U2002 ( .A(n69), .B(n1216), .C(n1215), .D(n66), .Z(n936) );
  COND2X1 U2003 ( .A(n69), .B(n1219), .C(n66), .D(n1218), .Z(n939) );
  CANR1XL U2004 ( .A(n278), .B(n287), .C(n279), .Z(n277) );
  CENX1 U2005 ( .A(n1715), .B(n152), .Z(n1280) );
  CENX1 U2006 ( .A(n1711), .B(n152), .Z(n1307) );
  CENX1 U2007 ( .A(n1698), .B(n152), .Z(n1400) );
  COND2X1 U2008 ( .A(n1175), .B(n1661), .C(n1176), .D(n91), .Z(n899) );
  CENX1 U2009 ( .A(a[16]), .B(n1734), .Z(n1445) );
  COND2XL U2010 ( .A(n85), .B(n1181), .C(n1657), .D(n1180), .Z(n903) );
  COND2XL U2011 ( .A(n85), .B(n1182), .C(n1181), .D(n1657), .Z(n904) );
  CNR2IX1 U2012 ( .B(n1691), .A(n1657), .Z(n916) );
  COND2XL U2013 ( .A(n85), .B(n1739), .C(n1657), .D(n1194), .Z(n851) );
  CENX1 U2014 ( .A(n1693), .B(n104), .Z(n1144) );
  COND2X1 U2015 ( .A(n36), .B(n1313), .C(n1312), .D(n1621), .Z(n1029) );
  CIVX1 U2016 ( .A(n1719), .Z(n1715) );
  COND2X1 U2017 ( .A(n53), .B(n1259), .C(n1624), .D(n1258), .Z(n977) );
  COND2XL U2018 ( .A(n61), .B(n1725), .C(n1251), .D(n58), .Z(n854) );
  COND2XL U2019 ( .A(n18), .B(n1659), .C(n1386), .D(n15), .Z(n859) );
  CENX1 U2020 ( .A(n1703), .B(n1684), .Z(n1374) );
  CENX1 U2021 ( .A(n1703), .B(n1685), .Z(n1372) );
  CENX1 U2022 ( .A(n1700), .B(b[24]), .Z(n1361) );
  CNR2XL U2023 ( .A(n294), .B(n291), .Z(n289) );
  CNR2X1 U2024 ( .A(n626), .B(n645), .Z(n263) );
  COND2XL U2025 ( .A(n53), .B(n1259), .C(n1624), .D(n1258), .Z(n1658) );
  CND2XL U2026 ( .A(n388), .B(n264), .Z(n175) );
  COND2XL U2027 ( .A(n18), .B(n1367), .C(n1366), .D(n15), .Z(n1081) );
  CND2IXL U2028 ( .B(n1691), .A(n1699), .Z(n1386) );
  CENX1 U2029 ( .A(n1699), .B(b[26]), .Z(n1359) );
  CIVX1 U2030 ( .A(n1713), .Z(n1710) );
  CENX1 U2031 ( .A(n1686), .B(n1731), .Z(n1195) );
  CIVXL U2032 ( .A(n12), .Z(n1659) );
  CFA1XL U2033 ( .A(n895), .B(n1105), .CI(n997), .CO(n523), .S(n524) );
  CIVX1 U2034 ( .A(n1713), .Z(n1711) );
  COND2XL U2035 ( .A(n18), .B(n1368), .C(n1367), .D(n15), .Z(n1082) );
  CENX1 U2036 ( .A(n1700), .B(n1686), .Z(n1370) );
  COND2XL U2037 ( .A(n44), .B(n1280), .C(n1279), .D(n42), .Z(n997) );
  COND2XL U2038 ( .A(n44), .B(n1279), .C(n1278), .D(n42), .Z(n996) );
  CND2IXL U2039 ( .B(n1691), .A(n1717), .Z(n1299) );
  CIVX2 U2040 ( .A(n1720), .Z(n1717) );
  CIVXL U2041 ( .A(n220), .Z(n222) );
  CIVX2 U2042 ( .A(n1728), .Z(n1727) );
  CNR2X1 U2043 ( .A(n280), .B(n285), .Z(n278) );
  CENX1 U2044 ( .A(n1680), .B(n1727), .Z(n1222) );
  COND2XL U2045 ( .A(n69), .B(n1728), .C(n1230), .D(n66), .Z(n853) );
  CENX1 U2046 ( .A(n1727), .B(n1681), .Z(n1221) );
  CENX1 U2047 ( .A(n1727), .B(n1677), .Z(n1225) );
  COND2XL U2048 ( .A(n44), .B(n1288), .C(n42), .D(n1287), .Z(n1005) );
  CENX1 U2049 ( .A(n1735), .B(a[20]), .Z(n1661) );
  COND2XL U2050 ( .A(n77), .B(n1205), .C(n1204), .D(n1557), .Z(n926) );
  CIVX2 U2051 ( .A(n1739), .Z(n1736) );
  CIVX1 U2052 ( .A(n1659), .Z(n1700) );
  CIVX1 U2053 ( .A(n1659), .Z(n1701) );
  CND2X1 U2054 ( .A(n534), .B(n557), .Z(n231) );
  CNR2X1 U2055 ( .A(n225), .B(n230), .Z(n219) );
  CND2X1 U2056 ( .A(n1640), .B(n1639), .Z(n236) );
  CND2XL U2057 ( .A(n1640), .B(n241), .Z(n172) );
  CNR2X1 U2058 ( .A(n236), .B(n252), .Z(n234) );
  CENX1 U2059 ( .A(n242), .B(n172), .Z(product[25]) );
  CND2XL U2060 ( .A(n1639), .B(n250), .Z(n173) );
  CND2XL U2061 ( .A(n606), .B(n608), .Z(n1673) );
  CND2X1 U2062 ( .A(n454), .B(n481), .Z(n210) );
  CANR1XL U2063 ( .A(n219), .B(n232), .C(n220), .Z(n218) );
  CANR1XL U2064 ( .A(n384), .B(n232), .C(n229), .Z(n227) );
  CND2XL U2065 ( .A(n384), .B(n231), .Z(n171) );
  CIVX1 U2066 ( .A(n231), .Z(n229) );
  CIVX1 U2067 ( .A(n230), .Z(n384) );
  CND2XL U2068 ( .A(n1049), .B(n939), .Z(n1662) );
  CND2XL U2069 ( .A(n1049), .B(n977), .Z(n1663) );
  CND2XL U2070 ( .A(n939), .B(n1658), .Z(n1664) );
  COND1XL U2071 ( .A(n294), .B(n307), .C(n295), .Z(n293) );
  CND2XL U2072 ( .A(n207), .B(n219), .Z(n205) );
  CEO3XL U2073 ( .A(n910), .B(n1050), .C(n958), .Z(n596) );
  CND2X1 U2074 ( .A(n910), .B(n1050), .Z(n1666) );
  CND2X1 U2075 ( .A(n910), .B(n958), .Z(n1667) );
  CND2XL U2076 ( .A(n600), .B(n615), .Z(n1669) );
  CND2XL U2077 ( .A(n600), .B(n596), .Z(n1670) );
  CND2XL U2078 ( .A(n615), .B(n596), .Z(n1671) );
  COND2XL U2079 ( .A(n27), .B(n1328), .C(n1327), .D(n1623), .Z(n1043) );
  COND2XL U2080 ( .A(n27), .B(n1329), .C(n1328), .D(n1623), .Z(n1044) );
  CIVX2 U2081 ( .A(n1734), .Z(n1733) );
  CND2XL U2082 ( .A(n606), .B(n627), .Z(n1672) );
  CND2XL U2083 ( .A(n627), .B(n608), .Z(n1674) );
  CND3XL U2084 ( .A(n1672), .B(n1673), .C(n1674), .Z(n603) );
  CND2X1 U2085 ( .A(n582), .B(n603), .Z(n250) );
  COND2XL U2086 ( .A(n77), .B(n1196), .C(n1557), .D(n1195), .Z(n917) );
  COND2XL U2087 ( .A(n1207), .B(n1557), .C(n1208), .D(n77), .Z(n929) );
  COND2XL U2088 ( .A(n77), .B(n1734), .C(n1557), .D(n1211), .Z(n852) );
  COND2XL U2089 ( .A(n77), .B(n1204), .C(n1557), .D(n1203), .Z(n925) );
  CND2IXL U2090 ( .B(n1691), .A(n1614), .Z(n1230) );
  COND2XL U2091 ( .A(n91), .B(n1168), .C(n1661), .D(n1167), .Z(n891) );
  COND2XL U2092 ( .A(n91), .B(n1169), .C(n1168), .D(n1661), .Z(n892) );
  COND2XL U2093 ( .A(n91), .B(n1170), .C(n1661), .D(n1169), .Z(n893) );
  COND2XL U2094 ( .A(n1177), .B(n1661), .C(n91), .D(n1178), .Z(n901) );
  COND2XL U2095 ( .A(n1171), .B(n1661), .C(n1172), .D(n91), .Z(n895) );
  COND2XL U2096 ( .A(n1171), .B(n91), .C(n1170), .D(n1661), .Z(n894) );
  CNR2IXL U2097 ( .B(n1691), .A(n1661), .Z(n902) );
  COND2XL U2098 ( .A(n1173), .B(n91), .C(n1172), .D(n1661), .Z(n896) );
  COND2XL U2099 ( .A(n1173), .B(n1661), .C(n1174), .D(n91), .Z(n897) );
  COND2XL U2100 ( .A(n1177), .B(n91), .C(n1176), .D(n1661), .Z(n900) );
  COND2XL U2101 ( .A(n91), .B(n1468), .C(n1661), .D(n1179), .Z(n850) );
  CND2IXL U2102 ( .B(n1691), .A(n1735), .Z(n1194) );
  CIVXL U2103 ( .A(n1705), .Z(n1699) );
  CIVXL U2104 ( .A(n1705), .Z(n1703) );
  CIVXL U2105 ( .A(n1705), .Z(n1704) );
  CIVXL U2106 ( .A(n1553), .Z(n1706) );
  CIVXL U2107 ( .A(n1553), .Z(n1708) );
  CIVXL U2108 ( .A(n1714), .Z(n1712) );
  CIVXL U2109 ( .A(n39), .Z(n1718) );
  CIVXL U2110 ( .A(n39), .Z(n1720) );
  CIVXL U2111 ( .A(n1739), .Z(n1737) );
  CIVX2 U2112 ( .A(n369), .Z(n407) );
  CIVX2 U2113 ( .A(n361), .Z(n405) );
  CIVX2 U2114 ( .A(n353), .Z(n403) );
  CIVX2 U2115 ( .A(n349), .Z(n402) );
  CIVX2 U2116 ( .A(n346), .Z(n401) );
  CIVX2 U2117 ( .A(n327), .Z(n398) );
  CIVX2 U2118 ( .A(n324), .Z(n397) );
  CIVX2 U2119 ( .A(n291), .Z(n392) );
  CIVX2 U2120 ( .A(n225), .Z(n383) );
  CIVX2 U2121 ( .A(n214), .Z(n382) );
  CIVX2 U2122 ( .A(n378), .Z(n376) );
  CIVX2 U2123 ( .A(n375), .Z(n373) );
  CIVX2 U2124 ( .A(n367), .Z(n365) );
  CIVX2 U2125 ( .A(n359), .Z(n357) );
  CIVX2 U2126 ( .A(n352), .Z(n351) );
  CIVX2 U2127 ( .A(n343), .Z(n342) );
  CIVX2 U2128 ( .A(n341), .Z(n339) );
  CIVX2 U2129 ( .A(n336), .Z(n334) );
  CIVX2 U2130 ( .A(n330), .Z(n329) );
  CIVX2 U2131 ( .A(n319), .Z(n317) );
  CIVX2 U2132 ( .A(n314), .Z(n312) );
  CIVX2 U2133 ( .A(n308), .Z(n307) );
  CIVX2 U2134 ( .A(n302), .Z(n304) );
  CIVX2 U2135 ( .A(n301), .Z(n394) );
  CIVX2 U2136 ( .A(n286), .Z(n284) );
  CIVX2 U2137 ( .A(n285), .Z(n391) );
  CIVX2 U2138 ( .A(n276), .Z(n274) );
  CIVX2 U2139 ( .A(n263), .Z(n388) );
  CIVX2 U2140 ( .A(n261), .Z(n259) );
  CIVX2 U2141 ( .A(n252), .Z(n254) );
  CIVX2 U2142 ( .A(n250), .Z(n248) );
  CIVX2 U2143 ( .A(n241), .Z(n239) );
  CIVX2 U2144 ( .A(n203), .Z(n201) );
  CIVX2 U2145 ( .A(n1687), .Z(n1468) );
  CIVX2 U2146 ( .A(n1688), .Z(n1467) );
  CIVX2 U2147 ( .A(n104), .Z(n1465) );
  CIVX2 U2148 ( .A(n113), .Z(n1463) );
endmodule


module calc_DW_mult_uns_14 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n3, n9, n12, n15, n18, n21, n27, n30, n33, n36, n39, n42, n44, n48,
         n50, n53, n55, n58, n61, n63, n66, n69, n71, n74, n77, n79, n82, n85,
         n87, n89, n91, n93, n95, n97, n99, n100, n102, n104, n105, n107, n109,
         n110, n112, n113, n114, n115, n116, n122, n124, n126, n128, n130,
         n132, n134, n136, n138, n140, n142, n144, n146, n148, n150, n151,
         n152, n153, n154, n155, n156, n157, n167, n168, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n198, n199, n205, n207, n208, n210, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n226, n227, n228, n229,
         n231, n234, n235, n236, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n248, n249, n250, n251, n252, n253, n257, n259, n260,
         n261, n262, n263, n264, n268, n270, n271, n272, n273, n275, n278,
         n279, n280, n281, n283, n285, n286, n288, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n301, n303, n304, n305, n306,
         n308, n311, n312, n313, n314, n316, n318, n319, n320, n321, n322,
         n323, n324, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n343, n345, n346, n348,
         n350, n351, n352, n354, n356, n357, n358, n359, n360, n362, n364,
         n365, n366, n367, n368, n370, n372, n373, n374, n375, n376, n378,
         n380, n381, n383, n387, n388, n389, n390, n391, n394, n397, n399,
         n401, n402, n403, n404, n410, n412, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1455, n1457, n1468, n1470, n1471, n1472, n1473,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720;
  assign n3 = a[1];
  assign n12 = a[3];
  assign n21 = a[5];
  assign n30 = a[7];
  assign n39 = a[9];
  assign n48 = a[11];
  assign n55 = a[13];
  assign n63 = a[15];
  assign n71 = a[17];
  assign n79 = a[19];
  assign n87 = a[21];
  assign n93 = a[23];
  assign n99 = a[25];
  assign n104 = a[27];
  assign n109 = a[29];
  assign n113 = a[31];
  assign n116 = b[0];
  assign n122 = b[2];
  assign n124 = b[3];
  assign n126 = b[4];
  assign n128 = b[5];
  assign n130 = b[6];
  assign n132 = b[7];
  assign n134 = b[8];
  assign n136 = b[9];
  assign n138 = b[10];
  assign n140 = b[11];
  assign n142 = b[12];
  assign n144 = b[13];
  assign n146 = b[14];
  assign n148 = b[15];
  assign n150 = b[16];
  assign n151 = b[17];
  assign n152 = b[18];
  assign n153 = b[19];
  assign n154 = b[20];
  assign n155 = b[21];
  assign n156 = b[22];
  assign n157 = b[23];

  COND1X1 U197 ( .A(n262), .B(n245), .C(n246), .Z(n244) );
  COND1X1 U304 ( .A(n328), .B(n322), .C(n323), .Z(n321) );
  CNR2X2 U307 ( .A(n767), .B(n778), .Z(n322) );
  CEO3X2 U412 ( .A(n444), .B(n423), .C(n442), .Z(n419) );
  CEO3X2 U413 ( .A(n425), .B(n424), .C(n446), .Z(n420) );
  CEO3X2 U414 ( .A(n428), .B(n427), .C(n426), .Z(n421) );
  CEO3X2 U416 ( .A(n456), .B(n429), .C(n454), .Z(n423) );
  CEO3X2 U417 ( .A(n956), .B(n1022), .C(n1076), .Z(n424) );
  CEO3X2 U418 ( .A(n938), .B(n998), .C(n1106), .Z(n425) );
  CEO3X2 U419 ( .A(n922), .B(n976), .C(n1048), .Z(n426) );
  CEO3X2 U420 ( .A(n868), .B(n896), .C(n866), .Z(n427) );
  CEO3X2 U421 ( .A(n878), .B(n850), .C(n908), .Z(n428) );
  CFA1X1 U424 ( .A(n439), .B(n462), .CI(n437), .CO(n432), .S(n433) );
  CFA1X1 U425 ( .A(n441), .B(n464), .CI(n466), .CO(n434), .S(n435) );
  CFA1X1 U426 ( .A(n468), .B(n443), .CI(n445), .CO(n436), .S(n437) );
  CFA1X1 U427 ( .A(n472), .B(n470), .CI(n447), .CO(n438), .S(n439) );
  CFA1X1 U428 ( .A(n451), .B(n449), .CI(n474), .CO(n440), .S(n441) );
  CFA1X1 U429 ( .A(n457), .B(n453), .CI(n455), .CO(n442), .S(n443) );
  CFA1X1 U430 ( .A(n480), .B(n476), .CI(n478), .CO(n444), .S(n445) );
  CFA1X1 U431 ( .A(n1049), .B(n482), .CI(n484), .CO(n446), .S(n447) );
  CFA1X1 U432 ( .A(n957), .B(n1077), .CI(n1023), .CO(n448), .S(n449) );
  CFA1X1 U433 ( .A(n939), .B(n1107), .CI(n977), .CO(n450), .S(n451) );
  CFA1X1 U435 ( .A(n909), .B(n869), .CI(n887), .CO(n454), .S(n455) );
  CFA1X1 U436 ( .A(n867), .B(n879), .CI(n873), .CO(n456), .S(n457) );
  CFA1X1 U437 ( .A(n463), .B(n461), .CI(n488), .CO(n458), .S(n459) );
  CFA1X1 U438 ( .A(n467), .B(n490), .CI(n465), .CO(n460), .S(n461) );
  CFA1X1 U439 ( .A(n469), .B(n492), .CI(n494), .CO(n462), .S(n463) );
  CFA1X1 U440 ( .A(n473), .B(n471), .CI(n496), .CO(n464), .S(n465) );
  CFA1X1 U441 ( .A(n475), .B(n498), .CI(n500), .CO(n466), .S(n467) );
  CFA1X1 U442 ( .A(n481), .B(n477), .CI(n479), .CO(n468), .S(n469) );
  CFA1X1 U443 ( .A(n504), .B(n483), .CI(n502), .CO(n470), .S(n471) );
  CFA1X1 U444 ( .A(n510), .B(n506), .CI(n508), .CO(n472), .S(n473) );
  CFA1X1 U445 ( .A(n1050), .B(n485), .CI(n1078), .CO(n474), .S(n475) );
  CFA1X1 U446 ( .A(n940), .B(n1108), .CI(n978), .CO(n476), .S(n477) );
  CFA1X1 U448 ( .A(n898), .B(n1000), .CI(n924), .CO(n480), .S(n481) );
  CFA1X1 U449 ( .A(n880), .B(n910), .CI(n851), .CO(n482), .S(n483) );
  CHA1X1 U450 ( .A(n874), .B(n888), .CO(n484), .S(n485) );
  CFA1X1 U451 ( .A(n491), .B(n489), .CI(n514), .CO(n486), .S(n487) );
  CFA1X1 U452 ( .A(n495), .B(n516), .CI(n493), .CO(n488), .S(n489) );
  CFA1X1 U453 ( .A(n497), .B(n518), .CI(n520), .CO(n490), .S(n491) );
  CFA1X1 U454 ( .A(n501), .B(n499), .CI(n522), .CO(n492), .S(n493) );
  CFA1X1 U455 ( .A(n524), .B(n503), .CI(n526), .CO(n494), .S(n495) );
  CFA1X1 U456 ( .A(n509), .B(n505), .CI(n507), .CO(n496), .S(n497) );
  CFA1X1 U457 ( .A(n530), .B(n511), .CI(n528), .CO(n498), .S(n499) );
  CFA1X1 U458 ( .A(n536), .B(n532), .CI(n534), .CO(n500), .S(n501) );
  CFA1X1 U460 ( .A(n959), .B(n1109), .CI(n1001), .CO(n504), .S(n505) );
  CFA1X1 U461 ( .A(n911), .B(n1025), .CI(n925), .CO(n506), .S(n507) );
  CFA1X1 U462 ( .A(n889), .B(n941), .CI(n899), .CO(n508), .S(n509) );
  CFA1X1 U463 ( .A(n871), .B(n881), .CI(n875), .CO(n510), .S(n511) );
  CFA1X1 U464 ( .A(n517), .B(n515), .CI(n540), .CO(n512), .S(n513) );
  CFA1X1 U465 ( .A(n521), .B(n542), .CI(n519), .CO(n514), .S(n515) );
  CFA1X1 U466 ( .A(n546), .B(n544), .CI(n523), .CO(n516), .S(n517) );
  CFA1X1 U467 ( .A(n527), .B(n525), .CI(n548), .CO(n518), .S(n519) );
  CFA1X1 U468 ( .A(n533), .B(n550), .CI(n529), .CO(n520), .S(n521) );
  CFA1X1 U469 ( .A(n535), .B(n531), .CI(n552), .CO(n522), .S(n523) );
  CFA1X1 U470 ( .A(n558), .B(n554), .CI(n556), .CO(n524), .S(n525) );
  CFA1X1 U471 ( .A(n1080), .B(n560), .CI(n537), .CO(n526), .S(n527) );
  CFA1X1 U472 ( .A(n980), .B(n1110), .CI(n1052), .CO(n528), .S(n529) );
  CFA1X1 U473 ( .A(n876), .B(n1002), .CI(n960), .CO(n530), .S(n531) );
  CFA1X1 U475 ( .A(n852), .B(n926), .CI(n900), .CO(n534), .S(n535) );
  CHA1X1 U476 ( .A(n882), .B(n890), .CO(n536), .S(n537) );
  CFA1X1 U478 ( .A(n568), .B(n566), .CI(n545), .CO(n540), .S(n541) );
  CFA1X1 U479 ( .A(n570), .B(n547), .CI(n549), .CO(n542), .S(n543) );
  CFA1X1 U480 ( .A(n574), .B(n551), .CI(n572), .CO(n544), .S(n545) );
  CFA1X1 U481 ( .A(n557), .B(n553), .CI(n555), .CO(n546), .S(n547) );
  CFA1X1 U482 ( .A(n576), .B(n559), .CI(n561), .CO(n548), .S(n549) );
  CFA1X1 U483 ( .A(n582), .B(n578), .CI(n580), .CO(n550), .S(n551) );
  CFA1X1 U484 ( .A(n1053), .B(n584), .CI(n1081), .CO(n552), .S(n553) );
  CFA1X1 U485 ( .A(n961), .B(n1111), .CI(n1599), .CO(n554), .S(n555) );
  CFA1X1 U486 ( .A(n913), .B(n1561), .CI(n943), .CO(n556), .S(n557) );
  CFA1X1 U487 ( .A(n901), .B(n1003), .CI(n927), .CO(n558), .S(n559) );
  CFA1X1 U488 ( .A(n877), .B(n891), .CI(n883), .CO(n560), .S(n561) );
  CFA1X1 U489 ( .A(n567), .B(n565), .CI(n588), .CO(n562), .S(n563) );
  CFA1X1 U490 ( .A(n592), .B(n590), .CI(n569), .CO(n564), .S(n565) );
  CFA1X1 U491 ( .A(n594), .B(n571), .CI(n573), .CO(n566), .S(n567) );
  CFA1X1 U492 ( .A(n598), .B(n575), .CI(n596), .CO(n568), .S(n569) );
  CFA1X1 U493 ( .A(n581), .B(n577), .CI(n579), .CO(n570), .S(n571) );
  CFA1X1 U494 ( .A(n602), .B(n583), .CI(n600), .CO(n572), .S(n573) );
  CFA1X1 U495 ( .A(n585), .B(n604), .CI(n606), .CO(n574), .S(n575) );
  CFA1X1 U496 ( .A(n1004), .B(n1112), .CI(n1082), .CO(n576), .S(n577) );
  CFA1X1 U497 ( .A(n928), .B(n1054), .CI(n982), .CO(n578), .S(n579) );
  CHA1X1 U500 ( .A(n853), .B(n902), .CO(n584), .S(n585) );
  CFA1X1 U501 ( .A(n591), .B(n589), .CI(n610), .CO(n586), .S(n587) );
  CFA1X1 U502 ( .A(n614), .B(n612), .CI(n593), .CO(n588), .S(n589) );
  CFA1X1 U503 ( .A(n616), .B(n595), .CI(n597), .CO(n590), .S(n591) );
  CFA1X1 U504 ( .A(n601), .B(n599), .CI(n618), .CO(n592), .S(n593) );
  CFA1X1 U505 ( .A(n605), .B(n620), .CI(n603), .CO(n594), .S(n595) );
  CFA1X1 U506 ( .A(n624), .B(n607), .CI(n622), .CO(n596), .S(n597) );
  CFA1X1 U507 ( .A(n1645), .B(n626), .CI(n628), .CO(n598), .S(n599) );
  CFA1X1 U508 ( .A(n963), .B(n1113), .CI(n1005), .CO(n600), .S(n601) );
  CFA1X1 U509 ( .A(n929), .B(n1055), .CI(n983), .CO(n602), .S(n603) );
  CFA1X1 U510 ( .A(n915), .B(n1560), .CI(n945), .CO(n604), .S(n605) );
  CFA1X1 U511 ( .A(n885), .B(n903), .CI(n893), .CO(n606), .S(n607) );
  CFA1X1 U512 ( .A(n613), .B(n611), .CI(n632), .CO(n608), .S(n609) );
  CFA1X1 U513 ( .A(n617), .B(n634), .CI(n615), .CO(n610), .S(n611) );
  CFA1X1 U514 ( .A(n638), .B(n636), .CI(n619), .CO(n612), .S(n613) );
  CFA1X1 U515 ( .A(n623), .B(n640), .CI(n621), .CO(n614), .S(n615) );
  CFA1X1 U516 ( .A(n642), .B(n625), .CI(n627), .CO(n616), .S(n617) );
  CFA1X1 U517 ( .A(n648), .B(n644), .CI(n646), .CO(n618), .S(n619) );
  CFA1X1 U518 ( .A(n1084), .B(n629), .CI(n1114), .CO(n620), .S(n621) );
  CFA1X1 U521 ( .A(n916), .B(n1030), .CI(n946), .CO(n626), .S(n627) );
  CHA1X1 U522 ( .A(n854), .B(n904), .CO(n628), .S(n629) );
  CFA1X1 U523 ( .A(n635), .B(n633), .CI(n652), .CO(n630), .S(n631) );
  CFA1X1 U524 ( .A(n639), .B(n654), .CI(n637), .CO(n632), .S(n633) );
  CFA1X1 U525 ( .A(n658), .B(n656), .CI(n641), .CO(n634), .S(n635) );
  CFA1X1 U526 ( .A(n645), .B(n643), .CI(n660), .CO(n636), .S(n637) );
  CFA1X1 U527 ( .A(n662), .B(n647), .CI(n649), .CO(n638), .S(n639) );
  CFA1X1 U528 ( .A(n668), .B(n664), .CI(n666), .CO(n640), .S(n641) );
  CFA1X1 U529 ( .A(n965), .B(n1085), .CI(n1031), .CO(n642), .S(n643) );
  CFA1X1 U530 ( .A(n947), .B(n1115), .CI(n1007), .CO(n644), .S(n645) );
  CFA1X1 U531 ( .A(n931), .B(n1057), .CI(n985), .CO(n646), .S(n647) );
  CFA1X1 U532 ( .A(n895), .B(n917), .CI(n905), .CO(n648), .S(n649) );
  CFA1X1 U533 ( .A(n655), .B(n653), .CI(n672), .CO(n650), .S(n651) );
  CFA1X1 U534 ( .A(n659), .B(n674), .CI(n657), .CO(n652), .S(n653) );
  CFA1X1 U535 ( .A(n678), .B(n676), .CI(n661), .CO(n654), .S(n655) );
  CFA1X1 U536 ( .A(n665), .B(n663), .CI(n680), .CO(n656), .S(n657) );
  CFA1X1 U538 ( .A(n1086), .B(n686), .CI(n669), .CO(n660), .S(n661) );
  CFA1X1 U539 ( .A(n986), .B(n1116), .CI(n1058), .CO(n662), .S(n663) );
  CFA1X1 U540 ( .A(n906), .B(n1008), .CI(n966), .CO(n664), .S(n665) );
  CFA1X1 U541 ( .A(n918), .B(n1032), .CI(n948), .CO(n666), .S(n667) );
  CHA1X1 U542 ( .A(n932), .B(n855), .CO(n668), .S(n669) );
  CFA1X1 U543 ( .A(n675), .B(n673), .CI(n690), .CO(n670), .S(n671) );
  CFA1X1 U544 ( .A(n679), .B(n692), .CI(n677), .CO(n672), .S(n673) );
  CFA1X1 U545 ( .A(n681), .B(n694), .CI(n696), .CO(n674), .S(n675) );
  CFA1X1 U546 ( .A(n687), .B(n683), .CI(n685), .CO(n676), .S(n677) );
  CFA1X1 U547 ( .A(n702), .B(n698), .CI(n700), .CO(n678), .S(n679) );
  CFA1X1 U548 ( .A(n1033), .B(n704), .CI(n1059), .CO(n680), .S(n681) );
  CFA1X1 U549 ( .A(n967), .B(n1087), .CI(n987), .CO(n682), .S(n683) );
  CFA1X1 U550 ( .A(n949), .B(n1117), .CI(n1009), .CO(n684), .S(n685) );
  CFA1X1 U552 ( .A(n693), .B(n691), .CI(n708), .CO(n688), .S(n689) );
  CFA1X1 U553 ( .A(n697), .B(n710), .CI(n695), .CO(n690), .S(n691) );
  CFA1X1 U554 ( .A(n699), .B(n712), .CI(n714), .CO(n692), .S(n693) );
  CFA1X1 U555 ( .A(n716), .B(n701), .CI(n703), .CO(n694), .S(n695) );
  CFA1X1 U556 ( .A(n705), .B(n718), .CI(n720), .CO(n696), .S(n697) );
  CFA1X1 U557 ( .A(n920), .B(n1088), .CI(n1034), .CO(n698), .S(n699) );
  CFA1X1 U558 ( .A(n950), .B(n1118), .CI(n1010), .CO(n700), .S(n701) );
  CHA1X1 U560 ( .A(n856), .B(n968), .CO(n704), .S(n705) );
  CFA1X1 U561 ( .A(n711), .B(n709), .CI(n724), .CO(n706), .S(n707) );
  CFA1X1 U562 ( .A(n715), .B(n726), .CI(n713), .CO(n708), .S(n709) );
  CFA1X1 U563 ( .A(n717), .B(n728), .CI(n730), .CO(n710), .S(n711) );
  CFA1X1 U564 ( .A(n732), .B(n719), .CI(n721), .CO(n712), .S(n713) );
  CFA1X1 U565 ( .A(n1061), .B(n734), .CI(n736), .CO(n714), .S(n715) );
  CFA1X1 U566 ( .A(n989), .B(n1089), .CI(n1035), .CO(n716), .S(n717) );
  CFA1X1 U567 ( .A(n969), .B(n1119), .CI(n1011), .CO(n718), .S(n719) );
  CFA1X1 U568 ( .A(n921), .B(n951), .CI(n935), .CO(n720), .S(n721) );
  CFA1X1 U569 ( .A(n727), .B(n725), .CI(n740), .CO(n722), .S(n723) );
  CFA1X1 U570 ( .A(n731), .B(n742), .CI(n729), .CO(n724), .S(n725) );
  CFA1X1 U571 ( .A(n735), .B(n744), .CI(n733), .CO(n726), .S(n727) );
  CFA1X1 U572 ( .A(n750), .B(n746), .CI(n748), .CO(n728), .S(n729) );
  CFA1X1 U573 ( .A(n1036), .B(n737), .CI(n1062), .CO(n730), .S(n731) );
  CFA1X1 U574 ( .A(n936), .B(n1557), .CI(n970), .CO(n732), .S(n733) );
  CFA1X1 U575 ( .A(n952), .B(n1120), .CI(n990), .CO(n734), .S(n735) );
  CHA1X1 U576 ( .A(n857), .B(n1012), .CO(n736), .S(n737) );
  CFA1X1 U577 ( .A(n743), .B(n741), .CI(n754), .CO(n738), .S(n739) );
  CFA1X1 U578 ( .A(n758), .B(n756), .CI(n745), .CO(n740), .S(n741) );
  CFA1X1 U579 ( .A(n751), .B(n747), .CI(n749), .CO(n742), .S(n743) );
  CFA1X1 U580 ( .A(n764), .B(n760), .CI(n762), .CO(n744), .S(n745) );
  CFA1X1 U581 ( .A(n1013), .B(n1091), .CI(n1063), .CO(n746), .S(n747) );
  CFA1X1 U582 ( .A(n991), .B(n1121), .CI(n1037), .CO(n748), .S(n749) );
  CFA1X1 U583 ( .A(n937), .B(n1595), .CI(n953), .CO(n750), .S(n751) );
  CFA1X1 U584 ( .A(n757), .B(n755), .CI(n768), .CO(n752), .S(n753) );
  CFA1X1 U585 ( .A(n772), .B(n759), .CI(n770), .CO(n754), .S(n755) );
  CFA1X1 U586 ( .A(n774), .B(n761), .CI(n763), .CO(n756), .S(n757) );
  CFA1X1 U587 ( .A(n1064), .B(n776), .CI(n765), .CO(n758), .S(n759) );
  CFA1X1 U588 ( .A(n972), .B(n1092), .CI(n1038), .CO(n760), .S(n761) );
  CFA1X1 U589 ( .A(n954), .B(n1122), .CI(n992), .CO(n762), .S(n763) );
  CHA1X1 U590 ( .A(n858), .B(n1014), .CO(n764), .S(n765) );
  CFA1X1 U591 ( .A(n771), .B(n769), .CI(n780), .CO(n766), .S(n767) );
  CFA1X1 U592 ( .A(n775), .B(n782), .CI(n773), .CO(n768), .S(n769) );
  CFA1X1 U593 ( .A(n786), .B(n777), .CI(n784), .CO(n770), .S(n771) );
  CFA1X1 U596 ( .A(n955), .B(n993), .CI(n973), .CO(n776), .S(n777) );
  CFA1X1 U597 ( .A(n783), .B(n781), .CI(n792), .CO(n778), .S(n779) );
  CFA1X1 U598 ( .A(n787), .B(n794), .CI(n785), .CO(n780), .S(n781) );
  CFA1X1 U599 ( .A(n789), .B(n796), .CI(n798), .CO(n782), .S(n783) );
  CFA1X1 U600 ( .A(n994), .B(n1094), .CI(n1066), .CO(n784), .S(n785) );
  CFA1X1 U601 ( .A(n974), .B(n1124), .CI(n1016), .CO(n786), .S(n787) );
  CHA1X1 U602 ( .A(n859), .B(n1040), .CO(n788), .S(n789) );
  CFA1X1 U603 ( .A(n802), .B(n793), .CI(n795), .CO(n790), .S(n791) );
  CFA1X1 U604 ( .A(n799), .B(n804), .CI(n797), .CO(n792), .S(n793) );
  CFA1X1 U605 ( .A(n1067), .B(n806), .CI(n808), .CO(n794), .S(n795) );
  CFA1X1 U606 ( .A(n1041), .B(n1125), .CI(n1095), .CO(n796), .S(n797) );
  CFA1X1 U607 ( .A(n975), .B(n1017), .CI(n995), .CO(n798), .S(n799) );
  CFA1X1 U608 ( .A(n805), .B(n803), .CI(n812), .CO(n800), .S(n801) );
  CFA1X1 U609 ( .A(n816), .B(n807), .CI(n814), .CO(n802), .S(n803) );
  CFA1X1 U610 ( .A(n1068), .B(n809), .CI(n1096), .CO(n804), .S(n805) );
  CFA1X1 U611 ( .A(n996), .B(n1126), .CI(n1597), .CO(n806), .S(n807) );
  CHA1X1 U612 ( .A(n860), .B(n1042), .CO(n808), .S(n809) );
  CFA1X1 U613 ( .A(n815), .B(n813), .CI(n820), .CO(n810), .S(n811) );
  CFA1X1 U614 ( .A(n824), .B(n817), .CI(n822), .CO(n812), .S(n813) );
  CFA1X1 U615 ( .A(n1069), .B(n1127), .CI(n1097), .CO(n814), .S(n815) );
  CFA1X1 U616 ( .A(n997), .B(n1043), .CI(n1019), .CO(n816), .S(n817) );
  CFA1X1 U617 ( .A(n823), .B(n821), .CI(n828), .CO(n818), .S(n819) );
  CFA1X1 U618 ( .A(n1044), .B(n830), .CI(n825), .CO(n820), .S(n821) );
  CFA1X1 U619 ( .A(n1020), .B(n1128), .CI(n1070), .CO(n822), .S(n823) );
  CHA1X1 U620 ( .A(n861), .B(n1098), .CO(n824), .S(n825) );
  CFA1X1 U621 ( .A(n834), .B(n829), .CI(n831), .CO(n826), .S(n827) );
  CFA1X1 U622 ( .A(n1099), .B(n836), .CI(n1129), .CO(n828), .S(n829) );
  CFA1X1 U624 ( .A(n837), .B(n835), .CI(n840), .CO(n832), .S(n833) );
  CFA1X1 U625 ( .A(n1046), .B(n1100), .CI(n1072), .CO(n834), .S(n835) );
  CHA1X1 U626 ( .A(n862), .B(n1130), .CO(n836), .S(n837) );
  CFA1X1 U627 ( .A(n1131), .B(n841), .CI(n844), .CO(n838), .S(n839) );
  CFA1X1 U629 ( .A(n1074), .B(n845), .CI(n1102), .CO(n842), .S(n843) );
  CHA1X1 U630 ( .A(n863), .B(n1132), .CO(n844), .S(n845) );
  CFA1X1 U631 ( .A(n1075), .B(n1133), .CI(n1103), .CO(n846), .S(n847) );
  CHA1X1 U632 ( .A(n864), .B(n1104), .CO(n848), .S(n849) );
  COND2X1 U633 ( .A(n115), .B(n1468), .C(n114), .D(n1139), .Z(n850) );
  COND2X1 U634 ( .A(n1138), .B(n115), .C(n114), .D(n1137), .Z(n866) );
  CND2IX1 U638 ( .B(n1675), .A(n113), .Z(n1139) );
  COND2X1 U639 ( .A(n112), .B(n1605), .C(n110), .D(n1144), .Z(n851) );
  COND2X1 U641 ( .A(n112), .B(n1142), .C(n110), .D(n1141), .Z(n869) );
  COND2X1 U642 ( .A(n1143), .B(n112), .C(n110), .D(n1142), .Z(n870) );
  COND2X1 U649 ( .A(n107), .B(n1470), .C(n105), .D(n1151), .Z(n852) );
  COND2X1 U651 ( .A(n107), .B(n1147), .C(n105), .D(n1146), .Z(n873) );
  COND2X1 U652 ( .A(n107), .B(n1148), .C(n105), .D(n1147), .Z(n874) );
  COND2X1 U653 ( .A(n107), .B(n1149), .C(n105), .D(n1148), .Z(n875) );
  COND2X1 U654 ( .A(n1150), .B(n107), .C(n105), .D(n1149), .Z(n876) );
  CND2IX1 U662 ( .B(n1675), .A(n104), .Z(n1151) );
  COND2X1 U667 ( .A(n102), .B(n1156), .C(n100), .D(n1155), .Z(n881) );
  COND2X1 U669 ( .A(n102), .B(n1158), .C(n100), .D(n1157), .Z(n883) );
  COND2X1 U670 ( .A(n1159), .B(n102), .C(n100), .D(n1158), .Z(n884) );
  CND2IX1 U680 ( .B(n1675), .A(n1673), .Z(n1160) );
  COND2X1 U681 ( .A(n97), .B(n1472), .C(n95), .D(n1171), .Z(n854) );
  COND2X1 U683 ( .A(n97), .B(n1163), .C(n1162), .D(n95), .Z(n887) );
  COND2X1 U687 ( .A(n97), .B(n1167), .C(n1166), .D(n95), .Z(n891) );
  COND2X1 U688 ( .A(n97), .B(n1168), .C(n1167), .D(n95), .Z(n892) );
  CND2IX1 U702 ( .B(n1675), .A(n1672), .Z(n1171) );
  COND2X1 U703 ( .A(n91), .B(n1473), .C(n89), .D(n1184), .Z(n855) );
  COND2X1 U708 ( .A(n91), .B(n1177), .C(n1176), .D(n89), .Z(n900) );
  COND2X1 U709 ( .A(n91), .B(n1178), .C(n1177), .D(n89), .Z(n901) );
  COND2X1 U710 ( .A(n91), .B(n1179), .C(n1178), .D(n89), .Z(n902) );
  COND2X1 U711 ( .A(n91), .B(n1180), .C(n1179), .D(n89), .Z(n903) );
  COND2X1 U712 ( .A(n91), .B(n1181), .C(n1180), .D(n89), .Z(n904) );
  COND2X1 U713 ( .A(n91), .B(n1182), .C(n1181), .D(n89), .Z(n905) );
  COND2X1 U714 ( .A(n1183), .B(n91), .C(n1182), .D(n89), .Z(n906) );
  CND2IX1 U728 ( .B(n1675), .A(n1621), .Z(n1184) );
  CND2IX1 U758 ( .B(n1675), .A(n1716), .Z(n1199) );
  COND2X1 U770 ( .A(n77), .B(n1211), .C(n1210), .D(n74), .Z(n932) );
  COND2X1 U798 ( .A(n69), .B(n1222), .C(n1221), .D(n66), .Z(n942) );
  COND2X1 U799 ( .A(n69), .B(n1223), .C(n1222), .D(n66), .Z(n943) );
  COND2X1 U800 ( .A(n69), .B(n1224), .C(n1223), .D(n66), .Z(n944) );
  COND2X1 U802 ( .A(n69), .B(n1226), .C(n1225), .D(n66), .Z(n946) );
  COND2X1 U803 ( .A(n69), .B(n1227), .C(n1226), .D(n66), .Z(n947) );
  COND2X1 U804 ( .A(n69), .B(n1228), .C(n1227), .D(n66), .Z(n948) );
  COND2X1 U805 ( .A(n69), .B(n1229), .C(n1228), .D(n66), .Z(n949) );
  COND2X1 U806 ( .A(n69), .B(n1230), .C(n1229), .D(n66), .Z(n950) );
  COND2X1 U807 ( .A(n69), .B(n1231), .C(n1230), .D(n66), .Z(n951) );
  COND2X1 U809 ( .A(n69), .B(n1233), .C(n1232), .D(n66), .Z(n953) );
  COND2X1 U810 ( .A(n69), .B(n1234), .C(n1233), .D(n66), .Z(n954) );
  COND2X1 U836 ( .A(n61), .B(n1241), .C(n1240), .D(n58), .Z(n960) );
  COND2X1 U837 ( .A(n61), .B(n1242), .C(n1241), .D(n58), .Z(n961) );
  COND2X1 U838 ( .A(n61), .B(n1243), .C(n1242), .D(n58), .Z(n962) );
  COND2X1 U839 ( .A(n61), .B(n1244), .C(n1243), .D(n58), .Z(n963) );
  COND2X1 U841 ( .A(n61), .B(n1246), .C(n1245), .D(n58), .Z(n965) );
  COND2X1 U842 ( .A(n61), .B(n1247), .C(n1246), .D(n58), .Z(n966) );
  COND2X1 U843 ( .A(n61), .B(n1248), .C(n1247), .D(n58), .Z(n967) );
  COND2X1 U844 ( .A(n61), .B(n1249), .C(n1248), .D(n58), .Z(n968) );
  COND2X1 U845 ( .A(n61), .B(n1250), .C(n1249), .D(n58), .Z(n969) );
  COND2X1 U848 ( .A(n61), .B(n1253), .C(n1252), .D(n58), .Z(n972) );
  COND2X1 U849 ( .A(n61), .B(n1254), .C(n1253), .D(n58), .Z(n973) );
  CND2IX1 U872 ( .B(n1675), .A(n1705), .Z(n1256) );
  COND2X1 U876 ( .A(n53), .B(n1260), .C(n1259), .D(n50), .Z(n978) );
  COND2X1 U880 ( .A(n53), .B(n1264), .C(n1263), .D(n50), .Z(n982) );
  COND2X1 U882 ( .A(n53), .B(n1266), .C(n1265), .D(n50), .Z(n984) );
  COND2X1 U883 ( .A(n53), .B(n1267), .C(n1266), .D(n50), .Z(n985) );
  COND2X1 U884 ( .A(n53), .B(n1268), .C(n1267), .D(n50), .Z(n986) );
  COND2X1 U885 ( .A(n53), .B(n1269), .C(n1268), .D(n50), .Z(n987) );
  COND2X1 U889 ( .A(n53), .B(n1273), .C(n1272), .D(n50), .Z(n991) );
  COND2X1 U890 ( .A(n53), .B(n1274), .C(n1273), .D(n50), .Z(n992) );
  COND2X1 U891 ( .A(n53), .B(n1275), .C(n1274), .D(n50), .Z(n993) );
  COND2X1 U893 ( .A(n53), .B(n1277), .C(n1276), .D(n50), .Z(n995) );
  COND2X1 U919 ( .A(n44), .B(n1700), .C(n1304), .D(n42), .Z(n861) );
  COND2X1 U920 ( .A(n44), .B(n1281), .C(n1280), .D(n42), .Z(n998) );
  COND2X1 U921 ( .A(n44), .B(n1282), .C(n1281), .D(n42), .Z(n999) );
  COND2X1 U922 ( .A(n44), .B(n1283), .C(n1282), .D(n42), .Z(n1000) );
  COND2X1 U923 ( .A(n44), .B(n1284), .C(n1283), .D(n42), .Z(n1001) );
  COND2X1 U924 ( .A(n44), .B(n1285), .C(n1284), .D(n42), .Z(n1002) );
  COND2X1 U925 ( .A(n44), .B(n1286), .C(n1285), .D(n42), .Z(n1003) );
  COND2X1 U926 ( .A(n44), .B(n1287), .C(n1286), .D(n42), .Z(n1004) );
  COND2X1 U928 ( .A(n44), .B(n1289), .C(n1288), .D(n42), .Z(n1006) );
  COND2X1 U929 ( .A(n44), .B(n1290), .C(n1289), .D(n42), .Z(n1007) );
  COND2X1 U930 ( .A(n44), .B(n1291), .C(n1290), .D(n42), .Z(n1008) );
  COND2X1 U931 ( .A(n44), .B(n1292), .C(n1291), .D(n42), .Z(n1009) );
  COND2X1 U932 ( .A(n44), .B(n1293), .C(n1292), .D(n42), .Z(n1010) );
  COND2X1 U933 ( .A(n44), .B(n1294), .C(n1293), .D(n42), .Z(n1011) );
  COND2X1 U934 ( .A(n44), .B(n1295), .C(n1294), .D(n42), .Z(n1012) );
  COND2X1 U935 ( .A(n44), .B(n1296), .C(n1295), .D(n42), .Z(n1013) );
  COND2X1 U936 ( .A(n44), .B(n1297), .C(n1296), .D(n42), .Z(n1014) );
  COND2X1 U937 ( .A(n44), .B(n1298), .C(n1297), .D(n42), .Z(n1015) );
  COND2X1 U938 ( .A(n44), .B(n1299), .C(n1298), .D(n42), .Z(n1016) );
  COND2X1 U939 ( .A(n44), .B(n1300), .C(n1299), .D(n42), .Z(n1017) );
  COND2X1 U941 ( .A(n44), .B(n1302), .C(n1301), .D(n42), .Z(n1019) );
  COND2X1 U942 ( .A(n44), .B(n1303), .C(n1302), .D(n42), .Z(n1020) );
  CND2IX1 U968 ( .B(n1675), .A(n1696), .Z(n1304) );
  COND2X1 U976 ( .A(n36), .B(n1312), .C(n1311), .D(n1655), .Z(n1028) );
  COND2X1 U978 ( .A(n36), .B(n1314), .C(n1313), .D(n1655), .Z(n1030) );
  COND2X1 U979 ( .A(n36), .B(n1315), .C(n1314), .D(n1655), .Z(n1031) );
  COND2X1 U980 ( .A(n36), .B(n1316), .C(n1315), .D(n1655), .Z(n1032) );
  COND2X1 U982 ( .A(n36), .B(n1318), .C(n1317), .D(n1655), .Z(n1034) );
  COND2X1 U985 ( .A(n36), .B(n1321), .C(n1320), .D(n1655), .Z(n1037) );
  COND2X1 U986 ( .A(n36), .B(n1322), .C(n1321), .D(n1655), .Z(n1038) );
  COND2X1 U988 ( .A(n36), .B(n1324), .C(n1323), .D(n1655), .Z(n1040) );
  COND2X1 U989 ( .A(n36), .B(n1325), .C(n1324), .D(n1655), .Z(n1041) );
  COND2X1 U990 ( .A(n36), .B(n1326), .C(n1325), .D(n1655), .Z(n1042) );
  COND2X1 U991 ( .A(n36), .B(n1327), .C(n1326), .D(n1655), .Z(n1043) );
  COND2X1 U1028 ( .A(n27), .B(n1337), .C(n1336), .D(n1559), .Z(n1052) );
  COND2X1 U1029 ( .A(n27), .B(n1338), .C(n1337), .D(n1559), .Z(n1053) );
  COND2X1 U1030 ( .A(n27), .B(n1339), .C(n1338), .D(n1559), .Z(n1054) );
  COND2X1 U1033 ( .A(n27), .B(n1342), .C(n1341), .D(n1559), .Z(n1057) );
  COND2X1 U1034 ( .A(n27), .B(n1343), .C(n1342), .D(n1559), .Z(n1058) );
  COND2X1 U1039 ( .A(n27), .B(n1348), .C(n1347), .D(n1559), .Z(n1063) );
  COND2X1 U1087 ( .A(n18), .B(n1367), .C(n1366), .D(n15), .Z(n1081) );
  COND2X1 U1088 ( .A(n18), .B(n1368), .C(n1367), .D(n15), .Z(n1082) );
  COND2X1 U1091 ( .A(n18), .B(n1371), .C(n1370), .D(n15), .Z(n1085) );
  COND2X1 U1093 ( .A(n18), .B(n1373), .C(n1372), .D(n15), .Z(n1087) );
  COND2X1 U1097 ( .A(n18), .B(n1377), .C(n1376), .D(n15), .Z(n1091) );
  COND2X1 U1098 ( .A(n18), .B(n1378), .C(n1377), .D(n15), .Z(n1092) );
  COND2X1 U1101 ( .A(n18), .B(n1381), .C(n1380), .D(n15), .Z(n1095) );
  COND2X1 U1109 ( .A(n18), .B(n1389), .C(n1388), .D(n15), .Z(n1103) );
  COND2X1 U1143 ( .A(n1576), .B(n1566), .C(n1676), .D(n1424), .Z(n865) );
  COND2X1 U1144 ( .A(n1576), .B(n1393), .C(n1676), .D(n1392), .Z(n1106) );
  COND2X1 U1145 ( .A(n1576), .B(n1394), .C(n1676), .D(n1393), .Z(n1107) );
  COND2X1 U1146 ( .A(n1576), .B(n1395), .C(n1676), .D(n1394), .Z(n1108) );
  COND2X1 U1147 ( .A(n1576), .B(n1396), .C(n1676), .D(n1395), .Z(n1109) );
  COND2X1 U1149 ( .A(n1576), .B(n1398), .C(n1676), .D(n1397), .Z(n1111) );
  COND2X1 U1150 ( .A(n1576), .B(n1399), .C(n1676), .D(n1398), .Z(n1112) );
  COND2X1 U1151 ( .A(n1654), .B(n1400), .C(n1676), .D(n1399), .Z(n1113) );
  COND2X1 U1152 ( .A(n1576), .B(n1401), .C(n1676), .D(n1400), .Z(n1114) );
  COND2X1 U1153 ( .A(n1654), .B(n1402), .C(n1676), .D(n1401), .Z(n1115) );
  COND2X1 U1154 ( .A(n1576), .B(n1403), .C(n1677), .D(n1402), .Z(n1116) );
  COND2X1 U1155 ( .A(n1654), .B(n1404), .C(n1677), .D(n1403), .Z(n1117) );
  COND2X1 U1156 ( .A(n1576), .B(n1405), .C(n1677), .D(n1404), .Z(n1118) );
  COND2X1 U1157 ( .A(n1654), .B(n1406), .C(n1677), .D(n1405), .Z(n1119) );
  COND2X1 U1158 ( .A(n1576), .B(n1407), .C(n1676), .D(n1406), .Z(n1120) );
  COND2X1 U1159 ( .A(n1654), .B(n1408), .C(n1676), .D(n1407), .Z(n1121) );
  COND2X1 U1160 ( .A(n1654), .B(n1409), .C(n1676), .D(n1408), .Z(n1122) );
  COND2X1 U1161 ( .A(n1576), .B(n1410), .C(n1676), .D(n1409), .Z(n1123) );
  COND2X1 U1162 ( .A(n1576), .B(n1411), .C(n1676), .D(n1410), .Z(n1124) );
  COND2X1 U1163 ( .A(n1576), .B(n1412), .C(n1676), .D(n1411), .Z(n1125) );
  COND2X1 U1164 ( .A(n1576), .B(n1413), .C(n1676), .D(n1412), .Z(n1126) );
  COND2X1 U1165 ( .A(n1576), .B(n1414), .C(n1676), .D(n1413), .Z(n1127) );
  COND2X1 U1166 ( .A(n1576), .B(n1415), .C(n1676), .D(n1414), .Z(n1128) );
  COND2X1 U1167 ( .A(n1576), .B(n1416), .C(n1676), .D(n1415), .Z(n1129) );
  COND2X1 U1168 ( .A(n1576), .B(n1417), .C(n1676), .D(n1416), .Z(n1130) );
  COND2X1 U1169 ( .A(n1576), .B(n1418), .C(n1676), .D(n1417), .Z(n1131) );
  COND2X1 U1170 ( .A(n1576), .B(n1419), .C(n1676), .D(n1418), .Z(n1132) );
  COND2X1 U1171 ( .A(n1576), .B(n1420), .C(n1676), .D(n1419), .Z(n1133) );
  COND2X1 U1172 ( .A(n1576), .B(n1421), .C(n1676), .D(n1420), .Z(n1134) );
  COND2X1 U1173 ( .A(n1576), .B(n1422), .C(n1676), .D(n1421), .Z(n1135) );
  COND2X1 U1174 ( .A(n1576), .B(n1423), .C(n1676), .D(n1422), .Z(n1136) );
  CND2IX1 U1208 ( .B(n1675), .A(n1567), .Z(n1424) );
  CEOX2 U1259 ( .A(a[12]), .B(n1705), .Z(n1452) );
  CIVX2 U1281 ( .A(n113), .Z(n1137) );
  CIVX2 U1282 ( .A(n1672), .Z(n1169) );
  CIVX2 U1283 ( .A(n1704), .Z(n1254) );
  CIVX2 U1284 ( .A(n1717), .Z(n1197) );
  CIVX2 U1285 ( .A(n1673), .Z(n1158) );
  CIVX2 U1286 ( .A(n104), .Z(n1149) );
  CIVX2 U1287 ( .A(n1617), .Z(n1302) );
  CIVX2 U1288 ( .A(n1621), .Z(n1182) );
  CIVX2 U1289 ( .A(n1683), .Z(n1389) );
  CIVX2 U1290 ( .A(n1713), .Z(n1214) );
  CIVX2 U1291 ( .A(n1563), .Z(n1329) );
  CIVX2 U1292 ( .A(n1708), .Z(n1233) );
  CIVX2 U1293 ( .A(n1679), .Z(n1422) );
  CIVX2 U1294 ( .A(n1701), .Z(n1277) );
  CENXL U1295 ( .A(1'b0), .B(n109), .Z(n1142) );
  CENXL U1296 ( .A(n1565), .B(1'b0), .Z(n1358) );
  COND2X1 U1297 ( .A(n61), .B(n1252), .C(n1251), .D(n58), .Z(n971) );
  CIVX3 U1298 ( .A(n1711), .Z(n1707) );
  CND2X2 U1299 ( .A(n1450), .B(n74), .Z(n77) );
  CNIVX4 U1300 ( .A(n116), .Z(n1675) );
  CENXL U1301 ( .A(n1696), .B(n155), .Z(n1282) );
  COND2XL U1302 ( .A(n36), .B(n1317), .C(n1316), .D(n1655), .Z(n1033) );
  CIVX1 U1303 ( .A(n1562), .Z(n1691) );
  CNR2IX1 U1304 ( .B(n1675), .A(n95), .Z(n895) );
  CNR2IX4 U1305 ( .B(n1675), .A(n89), .Z(n907) );
  CIVX1 U1306 ( .A(n262), .Z(n264) );
  COND1X1 U1307 ( .A(n214), .B(n242), .C(n215), .Z(n1573) );
  CNR2IX1 U1308 ( .B(n1675), .A(n66), .Z(n955) );
  CANR1X2 U1309 ( .A(n1635), .B(n321), .C(n316), .Z(n314) );
  CIVDX2 U1310 ( .A(n30), .Z0(n1562), .Z1(n1563) );
  CENXL U1311 ( .A(n1701), .B(n155), .Z(n1257) );
  CENX1 U1312 ( .A(n1692), .B(n155), .Z(n1309) );
  CNIVX4 U1313 ( .A(n93), .Z(n1672) );
  CENX1 U1314 ( .A(n1563), .B(n151), .Z(n1313) );
  CENX1 U1315 ( .A(n1565), .B(n151), .Z(n1342) );
  CENX1 U1316 ( .A(n1698), .B(n151), .Z(n1286) );
  CENX1 U1317 ( .A(n1680), .B(n151), .Z(n1373) );
  CENX1 U1318 ( .A(n1705), .B(n151), .Z(n1238) );
  CENX1 U1319 ( .A(n1565), .B(n1670), .Z(n1344) );
  CENXL U1320 ( .A(n1702), .B(n1670), .Z(n1263) );
  CNIVX2 U1321 ( .A(n148), .Z(n1670) );
  CENXL U1322 ( .A(n1659), .B(n104), .Z(n1146) );
  CENXL U1323 ( .A(n1679), .B(n1659), .Z(n1419) );
  CENXL U1324 ( .A(n1680), .B(n1659), .Z(n1386) );
  CENXL U1325 ( .A(n1659), .B(n1672), .Z(n1166) );
  CENXL U1326 ( .A(n1701), .B(n1659), .Z(n1274) );
  CNIVX1 U1327 ( .A(n1090), .Z(n1557) );
  COND2X1 U1328 ( .A(n85), .B(n1195), .C(n1194), .D(n82), .Z(n917) );
  CNIVX1 U1329 ( .A(n1628), .Z(n1558) );
  CNIVX2 U1330 ( .A(n1628), .Z(n1559) );
  CENX1 U1331 ( .A(n1681), .B(a[4]), .Z(n1628) );
  CANR1X2 U1332 ( .A(n229), .B(n216), .C(n217), .Z(n215) );
  CENXL U1333 ( .A(n1698), .B(n152), .Z(n1285) );
  CENXL U1334 ( .A(n1695), .B(n1670), .Z(n1315) );
  CND2X4 U1335 ( .A(n1455), .B(n1655), .Z(n36) );
  CFA1XL U1336 ( .A(n1039), .B(n788), .CI(n1093), .CO(n772), .S(n773) );
  CND3X1 U1337 ( .A(n1647), .B(n1648), .C(n1649), .Z(n658) );
  CND2XL U1338 ( .A(n667), .B(n682), .Z(n1648) );
  CNIVX1 U1339 ( .A(n1029), .Z(n1560) );
  CND3X1 U1340 ( .A(n1589), .B(n1590), .C(n1591), .Z(n582) );
  CNIVX1 U1341 ( .A(n1027), .Z(n1561) );
  CFA1XL U1342 ( .A(n1021), .B(n1071), .CI(n1045), .CO(n830), .S(n831) );
  CENXL U1343 ( .A(n1679), .B(n1665), .Z(n1413) );
  CENXL U1344 ( .A(n1622), .B(n1665), .Z(n1173) );
  CENXL U1345 ( .A(n1683), .B(n1665), .Z(n1380) );
  CENXL U1346 ( .A(n1713), .B(n1665), .Z(n1205) );
  CENXL U1347 ( .A(n1702), .B(n1665), .Z(n1268) );
  CENXL U1348 ( .A(n1702), .B(n151), .Z(n1261) );
  CENX1 U1349 ( .A(n1565), .B(n152), .Z(n1341) );
  CENXL U1350 ( .A(n1702), .B(n152), .Z(n1260) );
  CENXL U1351 ( .A(n1679), .B(n152), .Z(n1405) );
  CENXL U1352 ( .A(n1683), .B(n152), .Z(n1372) );
  CENXL U1353 ( .A(n1709), .B(n150), .Z(n1218) );
  CENXL U1354 ( .A(n1680), .B(n150), .Z(n1374) );
  CENXL U1355 ( .A(n1698), .B(n150), .Z(n1287) );
  CENXL U1356 ( .A(n1658), .B(n109), .Z(n1140) );
  CND2IX4 U1357 ( .B(n1626), .A(n42), .Z(n44) );
  COND2X2 U1358 ( .A(n44), .B(n1288), .C(n1287), .D(n42), .Z(n1005) );
  CIVX3 U1359 ( .A(n1646), .Z(n42) );
  CENX1 U1360 ( .A(n1657), .B(n1672), .Z(n1168) );
  CENX1 U1361 ( .A(n1717), .B(n1662), .Z(n1191) );
  CND2X1 U1362 ( .A(n1577), .B(n1578), .Z(n1060) );
  CND2X1 U1363 ( .A(n1579), .B(n1580), .Z(n1055) );
  CNIVX3 U1364 ( .A(n124), .Z(n1658) );
  CND2X1 U1365 ( .A(a[28]), .B(n1605), .Z(n1606) );
  CND2X1 U1366 ( .A(n1700), .B(n1618), .Z(n1620) );
  CENX1 U1367 ( .A(n1712), .B(n1660), .Z(n1210) );
  CENX1 U1368 ( .A(n1702), .B(n1666), .Z(n1267) );
  COR2X1 U1369 ( .A(n27), .B(n1340), .Z(n1579) );
  CENX1 U1370 ( .A(n1716), .B(n1660), .Z(n1193) );
  CENX1 U1371 ( .A(n1674), .B(n1673), .Z(n1159) );
  CENX1 U1372 ( .A(n1565), .B(n154), .Z(n1339) );
  CENX1 U1373 ( .A(n1701), .B(n1657), .Z(n1276) );
  CENX1 U1374 ( .A(n1701), .B(n1658), .Z(n1275) );
  CENX1 U1375 ( .A(n1679), .B(n1666), .Z(n1412) );
  CENX1 U1376 ( .A(n1697), .B(n1661), .Z(n1297) );
  CENX1 U1377 ( .A(n1701), .B(n1660), .Z(n1273) );
  CENX1 U1378 ( .A(n1704), .B(n1659), .Z(n1251) );
  CENX1 U1379 ( .A(n1567), .B(n151), .Z(n1406) );
  CENX1 U1380 ( .A(n1701), .B(n1661), .Z(n1272) );
  CENX1 U1381 ( .A(n1701), .B(n1663), .Z(n1270) );
  CENX1 U1382 ( .A(n1694), .B(n1666), .Z(n1319) );
  CENX1 U1383 ( .A(n1695), .B(n1668), .Z(n1317) );
  CENX1 U1384 ( .A(n1702), .B(n1664), .Z(n1269) );
  CENX1 U1385 ( .A(n1695), .B(n1669), .Z(n1316) );
  CENX1 U1386 ( .A(n1717), .B(n1658), .Z(n1195) );
  CENX1 U1387 ( .A(n1718), .B(n1664), .Z(n1189) );
  CNIVX1 U1388 ( .A(n138), .Z(n1665) );
  CENX1 U1389 ( .A(n1696), .B(n154), .Z(n1283) );
  CNIVX2 U1390 ( .A(n126), .Z(n1659) );
  CNIVX2 U1391 ( .A(n130), .Z(n1661) );
  CENX1 U1392 ( .A(n1679), .B(n1663), .Z(n1415) );
  CENX1 U1393 ( .A(n1679), .B(n1664), .Z(n1414) );
  CEOX1 U1394 ( .A(n1611), .B(n1616), .Z(n703) );
  CEOX1 U1395 ( .A(n1588), .B(n944), .Z(n583) );
  CEOX1 U1396 ( .A(n892), .B(n914), .Z(n1588) );
  CNIVX2 U1397 ( .A(n134), .Z(n1663) );
  CNIVX4 U1398 ( .A(n128), .Z(n1660) );
  CNIVX2 U1399 ( .A(n132), .Z(n1662) );
  CENX1 U1400 ( .A(n109), .B(a[30]), .Z(n114) );
  CNIVX2 U1401 ( .A(n140), .Z(n1666) );
  CENX1 U1402 ( .A(n1701), .B(n153), .Z(n1259) );
  CNIVX4 U1403 ( .A(n33), .Z(n1655) );
  CENX1 U1404 ( .A(n1689), .B(a[6]), .Z(n33) );
  CND2X2 U1405 ( .A(n1625), .B(n1558), .Z(n27) );
  CENX1 U1406 ( .A(n1679), .B(n1660), .Z(n1418) );
  CENX1 U1407 ( .A(n1679), .B(n1661), .Z(n1417) );
  CENX1 U1408 ( .A(n1679), .B(n1657), .Z(n1421) );
  CENX1 U1409 ( .A(n1679), .B(n1658), .Z(n1420) );
  CENX1 U1410 ( .A(n1679), .B(b[31]), .Z(n1392) );
  CEOX1 U1411 ( .A(n1600), .B(n433), .Z(n431) );
  CEOX1 U1412 ( .A(n435), .B(n460), .Z(n1600) );
  CND2X1 U1413 ( .A(n723), .B(n738), .Z(n303) );
  CND2X1 U1414 ( .A(n739), .B(n752), .Z(n306) );
  CNR2X2 U1415 ( .A(n707), .B(n722), .Z(n295) );
  CND2X1 U1416 ( .A(n689), .B(n706), .Z(n290) );
  CNR2X1 U1417 ( .A(n587), .B(n608), .Z(n249) );
  CND3XL U1418 ( .A(n1601), .B(n1602), .C(n1603), .Z(n430) );
  COND1XL U1419 ( .A(n223), .B(n231), .C(n226), .Z(n222) );
  CND2X1 U1420 ( .A(n459), .B(n486), .Z(n212) );
  CND2X1 U1421 ( .A(n431), .B(n458), .Z(n207) );
  CENX1 U1422 ( .A(n191), .B(n365), .Z(product[6]) );
  CENX1 U1423 ( .A(n1704), .B(n1658), .Z(n1252) );
  CENX1 U1424 ( .A(n1708), .B(n1657), .Z(n1232) );
  CENX1 U1425 ( .A(n1708), .B(n1658), .Z(n1231) );
  CIVX2 U1426 ( .A(n1711), .Z(n1708) );
  COND2X1 U1427 ( .A(n69), .B(n1232), .C(n1231), .D(n66), .Z(n952) );
  CIVDX1 U1428 ( .A(n21), .Z0(n1564), .Z1(n1565) );
  CIVX2 U1429 ( .A(n39), .Z(n1700) );
  CIVX2 U1430 ( .A(a[0]), .Z(n1677) );
  CIVX2 U1431 ( .A(a[0]), .Z(n1676) );
  CIVX2 U1432 ( .A(n71), .Z(n1715) );
  CIVX3 U1433 ( .A(n1715), .Z(n1712) );
  CIVDX2 U1434 ( .A(n3), .Z0(n1566), .Z1(n1567) );
  COR2X1 U1435 ( .A(n671), .B(n688), .Z(n1568) );
  COR2X1 U1436 ( .A(n631), .B(n650), .Z(n1569) );
  COR2X1 U1437 ( .A(n723), .B(n738), .Z(n1570) );
  CNIVX1 U1438 ( .A(n39), .Z(n1617) );
  COND2X1 U1439 ( .A(n85), .B(n1196), .C(n1195), .D(n82), .Z(n918) );
  COR2X1 U1440 ( .A(n431), .B(n458), .Z(n1571) );
  CAN2X1 U1441 ( .A(n1624), .B(n383), .Z(product[1]) );
  COND1X1 U1442 ( .A(n214), .B(n242), .C(n215), .Z(n213) );
  CANR1X1 U1443 ( .A(n1631), .B(n213), .C(n210), .Z(n208) );
  CENXL U1444 ( .A(n1574), .B(n220), .Z(product[28]) );
  CAN2XL U1445 ( .A(n387), .B(n219), .Z(n1574) );
  CENXL U1446 ( .A(n1565), .B(n155), .Z(n1338) );
  CENX2 U1447 ( .A(n1717), .B(n1657), .Z(n1196) );
  CENXL U1448 ( .A(n1575), .B(n199), .Z(product[31]) );
  CAN2X1 U1449 ( .A(n1639), .B(n198), .Z(n1575) );
  COND2XL U1450 ( .A(n36), .B(n1310), .C(n1309), .D(n1655), .Z(n1026) );
  COND2X1 U1451 ( .A(n97), .B(n1169), .C(n1168), .D(n95), .Z(n893) );
  CEOX2 U1452 ( .A(a[16]), .B(n1712), .Z(n1450) );
  CENXL U1453 ( .A(n1674), .B(n1702), .Z(n1278) );
  CND2IXL U1454 ( .B(n1675), .A(n1702), .Z(n1279) );
  CENX1 U1455 ( .A(n1708), .B(n1663), .Z(n1226) );
  CEOX1 U1456 ( .A(a[4]), .B(n1689), .Z(n1625) );
  COND2X1 U1457 ( .A(n27), .B(n1341), .C(n1340), .D(n1559), .Z(n1056) );
  COND2X1 U1458 ( .A(n85), .B(n1194), .C(n1193), .D(n82), .Z(n916) );
  COND2X1 U1459 ( .A(n77), .B(n1208), .C(n1207), .D(n74), .Z(n929) );
  CIVXL U1460 ( .A(n229), .Z(n231) );
  CNIVX4 U1461 ( .A(n9), .Z(n1576) );
  CND2IX2 U1462 ( .B(n1627), .A(n1676), .Z(n9) );
  COND2XL U1463 ( .A(n36), .B(n1306), .C(n1305), .D(n1655), .Z(n1022) );
  COND2XL U1464 ( .A(n36), .B(n1307), .C(n1306), .D(n1655), .Z(n1023) );
  COND2XL U1465 ( .A(n36), .B(n1328), .C(n1327), .D(n1655), .Z(n1044) );
  COND2XL U1466 ( .A(n36), .B(n1320), .C(n1319), .D(n1655), .Z(n1036) );
  COND2XL U1467 ( .A(n36), .B(n1330), .C(n1329), .D(n1655), .Z(n1046) );
  COND2XL U1468 ( .A(n36), .B(n1308), .C(n1307), .D(n1655), .Z(n1024) );
  COND2XL U1469 ( .A(n36), .B(n1323), .C(n1322), .D(n1655), .Z(n1039) );
  COND2XL U1470 ( .A(n36), .B(n1309), .C(n1308), .D(n1655), .Z(n1025) );
  COND2XL U1471 ( .A(n36), .B(n1329), .C(n1328), .D(n1655), .Z(n1045) );
  COND2XL U1472 ( .A(n36), .B(n1319), .C(n1318), .D(n1655), .Z(n1035) );
  CNR2IXL U1473 ( .B(n1675), .A(n1655), .Z(n1047) );
  COND2XL U1474 ( .A(n36), .B(n1311), .C(n1310), .D(n1655), .Z(n1027) );
  COND2XL U1475 ( .A(n36), .B(n1313), .C(n1312), .D(n1655), .Z(n1029) );
  CEOX2 U1476 ( .A(a[18]), .B(n1718), .Z(n1449) );
  CIVXL U1477 ( .A(n279), .Z(n278) );
  CIVX4 U1478 ( .A(n1685), .Z(n1681) );
  CFA1XL U1479 ( .A(n912), .B(n1026), .CI(n942), .CO(n532), .S(n533) );
  COND2X1 U1480 ( .A(n1170), .B(n97), .C(n95), .D(n1169), .Z(n894) );
  CENXL U1481 ( .A(n1674), .B(n1672), .Z(n1170) );
  CFA1X1 U1482 ( .A(n894), .B(n1006), .CI(n964), .CO(n624), .S(n625) );
  CENX1 U1483 ( .A(n1701), .B(n1668), .Z(n1265) );
  CANR1X1 U1484 ( .A(n228), .B(n241), .C(n229), .Z(n227) );
  CENXL U1485 ( .A(n1573), .B(n168), .Z(product[29]) );
  CFA1XL U1486 ( .A(n930), .B(n1056), .CI(n984), .CO(n622), .S(n623) );
  CANR1X1 U1487 ( .A(n390), .B(n241), .C(n238), .Z(n236) );
  CIVX2 U1488 ( .A(n242), .Z(n241) );
  CANR1X1 U1489 ( .A(n221), .B(n241), .C(n222), .Z(n220) );
  CEOX2 U1490 ( .A(a[6]), .B(n1563), .Z(n1455) );
  COND2X1 U1491 ( .A(n77), .B(n1212), .C(n1211), .D(n74), .Z(n933) );
  CIVDXL U1492 ( .A(n339), .Z0(n338) );
  CIVX2 U1493 ( .A(n1566), .Z(n1678) );
  CIVX2 U1494 ( .A(n63), .Z(n1711) );
  CENX1 U1495 ( .A(n1688), .B(n153), .Z(n1340) );
  COND2X1 U1496 ( .A(n69), .B(n1225), .C(n1224), .D(n66), .Z(n945) );
  COND1X1 U1497 ( .A(n226), .B(n218), .C(n219), .Z(n217) );
  COND2X1 U1498 ( .A(n1576), .B(n1397), .C(n1676), .D(n1396), .Z(n1110) );
  CND2X2 U1499 ( .A(n1446), .B(n100), .Z(n102) );
  CEOX1 U1500 ( .A(a[24]), .B(n1673), .Z(n1446) );
  COND2X1 U1501 ( .A(n102), .B(n1471), .C(n100), .D(n1160), .Z(n853) );
  CANR1X2 U1502 ( .A(n288), .B(n1568), .C(n283), .Z(n281) );
  CNR2IX1 U1503 ( .B(n1675), .A(n82), .Z(n921) );
  CANR1X2 U1504 ( .A(n257), .B(n391), .C(n248), .Z(n246) );
  CIVX1 U1505 ( .A(n250), .Z(n248) );
  CND2X2 U1506 ( .A(n391), .B(n1633), .Z(n245) );
  CENX4 U1507 ( .A(n1712), .B(a[18]), .Z(n82) );
  COND1X2 U1508 ( .A(n295), .B(n299), .C(n296), .Z(n294) );
  CNR2X1 U1509 ( .A(n295), .B(n298), .Z(n293) );
  CIVX4 U1510 ( .A(n1703), .Z(n1701) );
  COND1X2 U1511 ( .A(n330), .B(n313), .C(n314), .Z(n312) );
  COND2X1 U1512 ( .A(n18), .B(n1387), .C(n1386), .D(n15), .Z(n1101) );
  CIVX3 U1513 ( .A(n1566), .Z(n1679) );
  CND2X1 U1514 ( .A(n228), .B(n216), .Z(n214) );
  CNR2X1 U1515 ( .A(n234), .B(n239), .Z(n228) );
  CNR2X1 U1516 ( .A(n218), .B(n223), .Z(n216) );
  CENX2 U1517 ( .A(n1673), .B(a[26]), .Z(n105) );
  COR2XL U1518 ( .A(n1339), .B(n1559), .Z(n1580) );
  CND2X1 U1519 ( .A(n1570), .B(n399), .Z(n298) );
  CANR1X2 U1520 ( .A(n308), .B(n1570), .C(n301), .Z(n299) );
  CNR2X2 U1521 ( .A(n513), .B(n538), .Z(n223) );
  CIVX2 U1522 ( .A(n1720), .Z(n1718) );
  CIVX1 U1523 ( .A(n79), .Z(n1720) );
  CND2X2 U1524 ( .A(n1449), .B(n82), .Z(n85) );
  CANR1X1 U1525 ( .A(n1630), .B(n1573), .C(n1629), .Z(n199) );
  CENX4 U1526 ( .A(n1672), .B(a[24]), .Z(n100) );
  COND2X1 U1527 ( .A(n102), .B(n1155), .C(n100), .D(n1154), .Z(n880) );
  CNR2X2 U1528 ( .A(n1608), .B(n1609), .Z(n1610) );
  CIVX2 U1529 ( .A(n279), .Z(n1608) );
  COND1X2 U1530 ( .A(n240), .B(n234), .C(n235), .Z(n229) );
  CNR2X2 U1531 ( .A(n487), .B(n512), .Z(n218) );
  CEOX2 U1532 ( .A(a[10]), .B(n1702), .Z(n1453) );
  COR2XL U1533 ( .A(n27), .B(n1345), .Z(n1577) );
  COR2XL U1534 ( .A(n1344), .B(n1559), .Z(n1578) );
  CENXL U1535 ( .A(n1565), .B(n1669), .Z(n1345) );
  CEOX2 U1536 ( .A(n1060), .B(n1644), .Z(n1611) );
  CND2X1 U1537 ( .A(n1716), .B(a[20]), .Z(n1583) );
  CND2X1 U1538 ( .A(n1581), .B(n1582), .Z(n1584) );
  CND2X2 U1539 ( .A(n1583), .B(n1584), .Z(n89) );
  CIVX2 U1540 ( .A(n1716), .Z(n1581) );
  CIVX2 U1541 ( .A(a[20]), .Z(n1582) );
  COND2XL U1542 ( .A(n91), .B(n1174), .C(n1173), .D(n89), .Z(n897) );
  COND2XL U1543 ( .A(n91), .B(n1175), .C(n1174), .D(n89), .Z(n898) );
  COND2XL U1544 ( .A(n91), .B(n1176), .C(n1175), .D(n89), .Z(n899) );
  COND2XL U1545 ( .A(n91), .B(n1173), .C(n1172), .D(n89), .Z(n896) );
  CND2X1 U1546 ( .A(a[0]), .B(n1567), .Z(n1586) );
  CND2X2 U1547 ( .A(n1677), .B(n1585), .Z(n1587) );
  CND2X2 U1548 ( .A(n1586), .B(n1587), .Z(n1627) );
  CIVX2 U1549 ( .A(n1567), .Z(n1585) );
  CND2XL U1550 ( .A(n944), .B(n914), .Z(n1589) );
  CND2XL U1551 ( .A(n944), .B(n892), .Z(n1590) );
  CND2XL U1552 ( .A(n914), .B(n892), .Z(n1591) );
  COR2XL U1553 ( .A(n53), .B(n1262), .Z(n1592) );
  COR2XL U1554 ( .A(n1261), .B(n50), .Z(n1593) );
  CND2X1 U1555 ( .A(n1592), .B(n1593), .Z(n980) );
  CIVX1 U1556 ( .A(n971), .Z(n1594) );
  CIVX2 U1557 ( .A(n1594), .Z(n1595) );
  CNIVX1 U1558 ( .A(n87), .Z(n1621) );
  CNIVX1 U1559 ( .A(n87), .Z(n1622) );
  CNIVX4 U1560 ( .A(n87), .Z(n1671) );
  CFA1XL U1561 ( .A(n1047), .B(n1101), .CI(n1073), .CO(n840), .S(n841) );
  COND2XL U1562 ( .A(n102), .B(n1153), .C(n100), .D(n1152), .Z(n878) );
  COND2XL U1563 ( .A(n102), .B(n1154), .C(n100), .D(n1153), .Z(n879) );
  COND2XL U1564 ( .A(n102), .B(n1157), .C(n100), .D(n1156), .Z(n882) );
  CENXL U1565 ( .A(n1705), .B(n152), .Z(n1237) );
  CENXL U1566 ( .A(n1563), .B(n152), .Z(n1312) );
  COND2X1 U1567 ( .A(n85), .B(n1192), .C(n1191), .D(n82), .Z(n914) );
  CIVX4 U1568 ( .A(n1706), .Z(n1704) );
  CEOX2 U1569 ( .A(a[22]), .B(n1672), .Z(n1447) );
  CIVX1 U1570 ( .A(n1700), .Z(n1699) );
  CIVX1 U1571 ( .A(n1018), .Z(n1596) );
  CIVX2 U1572 ( .A(n1596), .Z(n1597) );
  CIVX2 U1573 ( .A(n1700), .Z(n1698) );
  CENXL U1574 ( .A(n1705), .B(n150), .Z(n1239) );
  CENXL U1575 ( .A(n1565), .B(n150), .Z(n1343) );
  CENXL U1576 ( .A(n1567), .B(n150), .Z(n1407) );
  CENXL U1577 ( .A(n1702), .B(n150), .Z(n1262) );
  CENXL U1578 ( .A(n1695), .B(n150), .Z(n1314) );
  CENXL U1579 ( .A(n1710), .B(n151), .Z(n1217) );
  CENXL U1580 ( .A(n1657), .B(n109), .Z(n1141) );
  CENXL U1581 ( .A(n1674), .B(n109), .Z(n1143) );
  CIVXL U1582 ( .A(n109), .Z(n1605) );
  CND2IXL U1583 ( .B(n1675), .A(n109), .Z(n1144) );
  CND2X1 U1584 ( .A(n1617), .B(a[10]), .Z(n1619) );
  CIVX2 U1585 ( .A(a[10]), .Z(n1618) );
  CIVX1 U1586 ( .A(n981), .Z(n1598) );
  CIVX2 U1587 ( .A(n1598), .Z(n1599) );
  CND2XL U1588 ( .A(n433), .B(n460), .Z(n1601) );
  CND2XL U1589 ( .A(n433), .B(n435), .Z(n1602) );
  CND2XL U1590 ( .A(n460), .B(n435), .Z(n1603) );
  CND2X1 U1591 ( .A(n1604), .B(n109), .Z(n1607) );
  CND2X2 U1592 ( .A(n1606), .B(n1607), .Z(n1444) );
  CIVXL U1593 ( .A(a[28]), .Z(n1604) );
  COND2XL U1594 ( .A(n112), .B(n1141), .C(n110), .D(n1140), .Z(n868) );
  CND2X2 U1595 ( .A(n1444), .B(n110), .Z(n112) );
  CNR2X2 U1596 ( .A(n1610), .B(n244), .Z(n242) );
  CIVX2 U1597 ( .A(n243), .Z(n1609) );
  CNR2X2 U1598 ( .A(n245), .B(n261), .Z(n243) );
  CND2XL U1599 ( .A(n988), .B(n1644), .Z(n1612) );
  CND2XL U1600 ( .A(n988), .B(n1060), .Z(n1613) );
  CND2XL U1601 ( .A(n1644), .B(n1060), .Z(n1614) );
  CND3X1 U1602 ( .A(n1612), .B(n1613), .C(n1614), .Z(n702) );
  CIVXL U1603 ( .A(n988), .Z(n1615) );
  CIVXL U1604 ( .A(n1615), .Z(n1616) );
  COND2XL U1605 ( .A(n53), .B(n1278), .C(n1277), .D(n50), .Z(n996) );
  COND2XL U1606 ( .A(n44), .B(n1301), .C(n1300), .D(n42), .Z(n1018) );
  CND2X4 U1607 ( .A(n1619), .B(n1620), .Z(n50) );
  COND2XL U1608 ( .A(n53), .B(n1270), .C(n1269), .D(n50), .Z(n988) );
  COND2XL U1609 ( .A(n53), .B(n1263), .C(n1262), .D(n50), .Z(n981) );
  COND2XL U1610 ( .A(n53), .B(n1272), .C(n1271), .D(n50), .Z(n990) );
  CND2X1 U1611 ( .A(n1568), .B(n1634), .Z(n280) );
  CNR2X1 U1612 ( .A(n322), .B(n327), .Z(n320) );
  CAN2XL U1613 ( .A(n1571), .B(n1631), .Z(n1630) );
  CENX1 U1614 ( .A(n1678), .B(n154), .Z(n1403) );
  CANR1X1 U1615 ( .A(n1638), .B(n357), .C(n354), .Z(n352) );
  CENXL U1616 ( .A(n1688), .B(n1664), .Z(n1350) );
  CENX1 U1617 ( .A(n1562), .B(a[8]), .Z(n1646) );
  CEOX1 U1618 ( .A(a[20]), .B(n1671), .Z(n1448) );
  CNR2X1 U1619 ( .A(n563), .B(n586), .Z(n239) );
  CND2X2 U1620 ( .A(n1569), .B(n394), .Z(n261) );
  CND2X1 U1621 ( .A(n801), .B(n810), .Z(n337) );
  COR2X1 U1622 ( .A(n819), .B(n826), .Z(n1636) );
  CANR1XL U1623 ( .A(n381), .B(n1643), .C(n378), .Z(n376) );
  CND2XL U1624 ( .A(n412), .B(n375), .Z(n194) );
  CND2XL U1625 ( .A(n410), .B(n367), .Z(n192) );
  CEO3X1 U1626 ( .A(n452), .B(n450), .C(n448), .Z(n422) );
  CENX1 U1627 ( .A(n1692), .B(n1662), .Z(n1323) );
  CENX1 U1628 ( .A(n1697), .B(n1662), .Z(n1296) );
  CENX1 U1629 ( .A(n1567), .B(n1669), .Z(n1409) );
  CNR2IX1 U1630 ( .B(n1675), .A(n110), .Z(n871) );
  CENX1 U1631 ( .A(n1565), .B(n1660), .Z(n1354) );
  CENX1 U1632 ( .A(n1701), .B(n1662), .Z(n1271) );
  CIVX2 U1633 ( .A(n1719), .Z(n1716) );
  CENX1 U1634 ( .A(a[8]), .B(n1699), .Z(n1626) );
  CENX1 U1635 ( .A(n1680), .B(b[24]), .Z(n1366) );
  CENX1 U1636 ( .A(n1684), .B(b[25]), .Z(n1365) );
  CENX1 U1637 ( .A(n1686), .B(b[24]), .Z(n1335) );
  CND2XL U1638 ( .A(n389), .B(n235), .Z(n171) );
  CEOXL U1639 ( .A(n227), .B(n170), .Z(product[27]) );
  CNR2IXL U1640 ( .B(n228), .A(n223), .Z(n221) );
  CND2XL U1641 ( .A(n1635), .B(n318), .Z(n182) );
  CEOXL U1642 ( .A(n182), .B(n319), .Z(product[15]) );
  CEOXL U1643 ( .A(n297), .B(n1623), .Z(product[18]) );
  CAN2XL U1644 ( .A(n397), .B(n296), .Z(n1623) );
  CND2XL U1645 ( .A(n320), .B(n1635), .Z(n313) );
  CIVX1 U1646 ( .A(n318), .Z(n316) );
  CIVX1 U1647 ( .A(n285), .Z(n283) );
  CEOXL U1648 ( .A(n177), .B(n286), .Z(product[20]) );
  CEOXL U1649 ( .A(n176), .B(n278), .Z(product[21]) );
  CEOXL U1650 ( .A(n183), .B(n324), .Z(product[14]) );
  CND2XL U1651 ( .A(n401), .B(n323), .Z(n183) );
  CEOXL U1652 ( .A(n181), .B(n311), .Z(product[16]) );
  CANR1X1 U1653 ( .A(n331), .B(n339), .C(n332), .Z(n330) );
  CNR2XL U1654 ( .A(n333), .B(n336), .Z(n331) );
  CND2XL U1655 ( .A(n1637), .B(n345), .Z(n187) );
  CND2XL U1656 ( .A(n1636), .B(n350), .Z(n188) );
  CND2XL U1657 ( .A(n402), .B(n328), .Z(n184) );
  CND2XL U1658 ( .A(n430), .B(n415), .Z(n198) );
  CND2XL U1659 ( .A(n1638), .B(n356), .Z(n189) );
  CND2IXL U1660 ( .B(n358), .A(n359), .Z(n190) );
  CND2XL U1661 ( .A(n1642), .B(n364), .Z(n191) );
  CND2XL U1662 ( .A(n791), .B(n800), .Z(n334) );
  CANR1X1 U1663 ( .A(n365), .B(n1642), .C(n362), .Z(n360) );
  CND2XL U1664 ( .A(n1643), .B(n380), .Z(n195) );
  CND2XL U1665 ( .A(n1640), .B(n372), .Z(n193) );
  CEOXL U1666 ( .A(n376), .B(n194), .Z(product[3]) );
  CEOXL U1667 ( .A(n368), .B(n192), .Z(product[5]) );
  CND2XL U1668 ( .A(n843), .B(n846), .Z(n367) );
  CND2XL U1669 ( .A(n849), .B(n1134), .Z(n375) );
  CEO3X1 U1670 ( .A(n434), .B(n416), .C(n432), .Z(n415) );
  CEO3X1 U1671 ( .A(n436), .B(n418), .C(n417), .Z(n416) );
  CEO3X1 U1672 ( .A(n422), .B(n421), .C(n440), .Z(n418) );
  CEO3X1 U1673 ( .A(n420), .B(n438), .C(n419), .Z(n417) );
  COR2XL U1674 ( .A(n1136), .B(n865), .Z(n1624) );
  CNR2IXL U1675 ( .B(n1675), .A(n100), .Z(n885) );
  CNR2IXL U1676 ( .B(n1675), .A(n105), .Z(n877) );
  CIVXL U1677 ( .A(n1711), .Z(n1709) );
  CNR2IXL U1678 ( .B(n1675), .A(n42), .Z(n1021) );
  COND2XL U1679 ( .A(n107), .B(n1146), .C(n105), .D(n1145), .Z(n872) );
  CNR2IXL U1680 ( .B(n1675), .A(n1676), .Z(product[0]) );
  CENX2 U1681 ( .A(n1671), .B(a[22]), .Z(n95) );
  CND2X2 U1682 ( .A(n95), .B(n1447), .Z(n97) );
  CENXL U1683 ( .A(n1705), .B(n153), .Z(n1236) );
  CEOXL U1684 ( .A(a[26]), .B(n104), .Z(n1445) );
  CNIVX4 U1685 ( .A(n122), .Z(n1657) );
  CENXL U1686 ( .A(n1701), .B(n154), .Z(n1258) );
  CND2XL U1687 ( .A(n1443), .B(n114), .Z(n115) );
  CIVX2 U1688 ( .A(n48), .Z(n1703) );
  CIVX2 U1689 ( .A(n55), .Z(n1706) );
  CND2XL U1690 ( .A(n1571), .B(n207), .Z(n167) );
  CENX1 U1691 ( .A(n241), .B(n172), .Z(product[25]) );
  CND2XL U1692 ( .A(n1631), .B(n212), .Z(n168) );
  CND2XL U1693 ( .A(n388), .B(n226), .Z(n170) );
  CAOR1X1 U1694 ( .A(n210), .B(n1571), .C(n205), .Z(n1629) );
  CNR2X1 U1695 ( .A(n539), .B(n562), .Z(n234) );
  CENX1 U1696 ( .A(n260), .B(n174), .Z(product[23]) );
  CND2X1 U1697 ( .A(n1633), .B(n259), .Z(n174) );
  CANR1XL U1698 ( .A(n1633), .B(n264), .C(n257), .Z(n253) );
  CENX1 U1699 ( .A(n291), .B(n178), .Z(product[19]) );
  CND2XL U1700 ( .A(n1634), .B(n290), .Z(n178) );
  CENX1 U1701 ( .A(n271), .B(n175), .Z(product[22]) );
  COND1XL U1702 ( .A(n272), .B(n278), .C(n273), .Z(n271) );
  CENX1 U1703 ( .A(n251), .B(n173), .Z(product[24]) );
  COND1XL U1704 ( .A(n252), .B(n278), .C(n253), .Z(n251) );
  CND2X1 U1705 ( .A(n263), .B(n1633), .Z(n252) );
  CENX1 U1706 ( .A(n304), .B(n180), .Z(product[17]) );
  CND2XL U1707 ( .A(n1570), .B(n303), .Z(n180) );
  COND1XL U1708 ( .A(n305), .B(n311), .C(n306), .Z(n304) );
  CND2XL U1709 ( .A(n1568), .B(n285), .Z(n177) );
  CANR1XL U1710 ( .A(n1634), .B(n291), .C(n288), .Z(n286) );
  CANR1XL U1711 ( .A(n402), .B(n329), .C(n326), .Z(n324) );
  CND2XL U1712 ( .A(n399), .B(n306), .Z(n181) );
  COR2X1 U1713 ( .A(n459), .B(n486), .Z(n1631) );
  CND2X1 U1714 ( .A(n563), .B(n586), .Z(n240) );
  CND2X1 U1715 ( .A(n587), .B(n608), .Z(n250) );
  COND1XL U1716 ( .A(n337), .B(n333), .C(n334), .Z(n332) );
  COND1XL U1717 ( .A(n352), .B(n340), .C(n341), .Z(n339) );
  CND2X1 U1718 ( .A(n1637), .B(n1636), .Z(n340) );
  CANR1XL U1719 ( .A(n348), .B(n1637), .C(n343), .Z(n341) );
  CENX1 U1720 ( .A(n1632), .B(n541), .Z(n539) );
  CENX1 U1721 ( .A(n543), .B(n564), .Z(n1632) );
  CND3XL U1722 ( .A(n1651), .B(n1652), .C(n1653), .Z(n538) );
  CENX1 U1723 ( .A(n188), .B(n351), .Z(product[9]) );
  CENX1 U1724 ( .A(n335), .B(n185), .Z(product[12]) );
  CND2X1 U1725 ( .A(n403), .B(n334), .Z(n185) );
  COND1XL U1726 ( .A(n336), .B(n338), .C(n337), .Z(n335) );
  CENX1 U1727 ( .A(n329), .B(n184), .Z(product[13]) );
  CNR2X1 U1728 ( .A(n739), .B(n752), .Z(n305) );
  COR2X1 U1729 ( .A(n609), .B(n630), .Z(n1633) );
  CEOX1 U1730 ( .A(n346), .B(n187), .Z(product[10]) );
  CANR1XL U1731 ( .A(n1636), .B(n351), .C(n348), .Z(n346) );
  CEOX1 U1732 ( .A(n186), .B(n338), .Z(product[11]) );
  CND2X1 U1733 ( .A(n404), .B(n337), .Z(n186) );
  COR2X1 U1734 ( .A(n689), .B(n706), .Z(n1634) );
  COR2X1 U1735 ( .A(n753), .B(n766), .Z(n1635) );
  CND2X1 U1736 ( .A(n671), .B(n688), .Z(n285) );
  CND2X1 U1737 ( .A(n609), .B(n630), .Z(n259) );
  CND2X1 U1738 ( .A(n753), .B(n766), .Z(n318) );
  CND2X1 U1739 ( .A(n707), .B(n722), .Z(n296) );
  CND2X1 U1740 ( .A(n767), .B(n778), .Z(n323) );
  CND2X1 U1741 ( .A(n651), .B(n670), .Z(n273) );
  CND2X1 U1742 ( .A(n631), .B(n650), .Z(n270) );
  COND1XL U1743 ( .A(n376), .B(n374), .C(n375), .Z(n373) );
  COND1XL U1744 ( .A(n358), .B(n360), .C(n359), .Z(n357) );
  COND1XL U1745 ( .A(n368), .B(n366), .C(n367), .Z(n365) );
  CANR1XL U1746 ( .A(n373), .B(n1640), .C(n370), .Z(n368) );
  CNR2X1 U1747 ( .A(n801), .B(n810), .Z(n336) );
  CNR2X1 U1748 ( .A(n791), .B(n800), .Z(n333) );
  CNR2X1 U1749 ( .A(n779), .B(n790), .Z(n327) );
  COR2X1 U1750 ( .A(n811), .B(n818), .Z(n1637) );
  CND2X1 U1751 ( .A(n779), .B(n790), .Z(n328) );
  CND2X1 U1752 ( .A(n819), .B(n826), .Z(n350) );
  CND2X1 U1753 ( .A(n827), .B(n832), .Z(n356) );
  CND2X1 U1754 ( .A(n811), .B(n818), .Z(n345) );
  COR2X1 U1755 ( .A(n827), .B(n832), .Z(n1638) );
  COR2X1 U1756 ( .A(n430), .B(n415), .Z(n1639) );
  CENX1 U1757 ( .A(n189), .B(n1650), .Z(product[8]) );
  CENX1 U1758 ( .A(n193), .B(n373), .Z(product[4]) );
  CENX1 U1759 ( .A(n195), .B(n381), .Z(product[2]) );
  CNR2X1 U1760 ( .A(n843), .B(n846), .Z(n366) );
  CNR2X1 U1761 ( .A(n833), .B(n838), .Z(n358) );
  CNR2X1 U1762 ( .A(n849), .B(n1134), .Z(n374) );
  COR2X1 U1763 ( .A(n847), .B(n848), .Z(n1640) );
  CENX1 U1764 ( .A(n1641), .B(n667), .Z(n659) );
  CENX1 U1765 ( .A(n682), .B(n684), .Z(n1641) );
  CND2X1 U1766 ( .A(n1136), .B(n865), .Z(n383) );
  CND2X1 U1767 ( .A(n1135), .B(n1105), .Z(n380) );
  CND2X1 U1768 ( .A(n847), .B(n848), .Z(n372) );
  CND2X1 U1769 ( .A(n839), .B(n842), .Z(n364) );
  COR2X1 U1770 ( .A(n839), .B(n842), .Z(n1642) );
  CND2X1 U1771 ( .A(n833), .B(n838), .Z(n359) );
  COR2X1 U1772 ( .A(n1135), .B(n1105), .Z(n1643) );
  CENX1 U1773 ( .A(n1672), .B(n1664), .Z(n1161) );
  CENX1 U1774 ( .A(n1717), .B(n1668), .Z(n1185) );
  CENX1 U1775 ( .A(n1563), .B(n1663), .Z(n1322) );
  CENX1 U1776 ( .A(n1707), .B(n1660), .Z(n1229) );
  CENX1 U1777 ( .A(n1707), .B(n1661), .Z(n1228) );
  CENX1 U1778 ( .A(n1693), .B(n1660), .Z(n1325) );
  CENX1 U1779 ( .A(n1692), .B(n1661), .Z(n1324) );
  CENX1 U1780 ( .A(n1694), .B(n1667), .Z(n1318) );
  CENX1 U1781 ( .A(n1707), .B(n1659), .Z(n1230) );
  CENX1 U1782 ( .A(n1693), .B(n1659), .Z(n1326) );
  CENX1 U1783 ( .A(n1713), .B(n1664), .Z(n1206) );
  CENX1 U1784 ( .A(n1708), .B(n1662), .Z(n1227) );
  CENX1 U1785 ( .A(n1693), .B(n1657), .Z(n1328) );
  CENX1 U1786 ( .A(n1697), .B(n1659), .Z(n1299) );
  CENX1 U1787 ( .A(n1694), .B(n1664), .Z(n1321) );
  CENX1 U1788 ( .A(n1710), .B(n1666), .Z(n1223) );
  CENX1 U1789 ( .A(n1674), .B(n1567), .Z(n1423) );
  CIVX2 U1790 ( .A(n1703), .Z(n1702) );
  CENX1 U1791 ( .A(n1712), .B(n1661), .Z(n1209) );
  CENX1 U1792 ( .A(n1714), .B(n1666), .Z(n1204) );
  CENX1 U1793 ( .A(n1713), .B(n1657), .Z(n1213) );
  CENX1 U1794 ( .A(n1707), .B(n1664), .Z(n1225) );
  CENX1 U1795 ( .A(n1682), .B(n1657), .Z(n1388) );
  CENX1 U1796 ( .A(n1622), .B(n1666), .Z(n1172) );
  CENX1 U1797 ( .A(n1713), .B(n1663), .Z(n1207) );
  CENX1 U1798 ( .A(n1710), .B(n1665), .Z(n1224) );
  CENX1 U1799 ( .A(n1712), .B(n1659), .Z(n1211) );
  CENX1 U1800 ( .A(n1687), .B(n1659), .Z(n1355) );
  CIVX2 U1801 ( .A(n1706), .Z(n1705) );
  CENX1 U1802 ( .A(n1714), .B(n1670), .Z(n1200) );
  CENX1 U1803 ( .A(n1675), .B(n1710), .Z(n1234) );
  CENX1 U1804 ( .A(n1674), .B(n1563), .Z(n1330) );
  CENX1 U1805 ( .A(n1682), .B(n1666), .Z(n1379) );
  CENX1 U1806 ( .A(n1690), .B(n1663), .Z(n1351) );
  CENX1 U1807 ( .A(n1718), .B(n1665), .Z(n1188) );
  CENX1 U1808 ( .A(n1718), .B(n1666), .Z(n1187) );
  CENX1 U1809 ( .A(n1714), .B(n1668), .Z(n1202) );
  CENX1 U1810 ( .A(n1714), .B(n1669), .Z(n1201) );
  CENX1 U1811 ( .A(n1717), .B(n1667), .Z(n1186) );
  CENX1 U1812 ( .A(n1710), .B(n1670), .Z(n1219) );
  CENX1 U1813 ( .A(n1718), .B(n1663), .Z(n1190) );
  CENX1 U1814 ( .A(n1713), .B(n1658), .Z(n1212) );
  CENX1 U1815 ( .A(n1683), .B(n1660), .Z(n1385) );
  CENX1 U1816 ( .A(n1688), .B(n1662), .Z(n1352) );
  CENX1 U1817 ( .A(n1684), .B(n1658), .Z(n1387) );
  CENX1 U1818 ( .A(n1662), .B(n1673), .Z(n1152) );
  CNR2IXL U1819 ( .B(n1675), .A(n15), .Z(n1105) );
  CENX1 U1820 ( .A(n1698), .B(n1664), .Z(n1294) );
  CENX1 U1821 ( .A(n1698), .B(n1663), .Z(n1295) );
  CENX1 U1822 ( .A(n1702), .B(n1667), .Z(n1266) );
  CENX1 U1823 ( .A(n1622), .B(n1657), .Z(n1181) );
  CENX1 U1824 ( .A(n1622), .B(n1662), .Z(n1176) );
  CENX1 U1825 ( .A(n1621), .B(n1661), .Z(n1177) );
  CENX1 U1826 ( .A(n1621), .B(n1664), .Z(n1174) );
  CENX1 U1827 ( .A(n1704), .B(n1662), .Z(n1248) );
  CENX1 U1828 ( .A(n1704), .B(n1657), .Z(n1253) );
  CENX1 U1829 ( .A(n1704), .B(n1663), .Z(n1247) );
  CENX1 U1830 ( .A(n1704), .B(n1661), .Z(n1249) );
  CENX1 U1831 ( .A(n1682), .B(n1668), .Z(n1377) );
  CENX1 U1832 ( .A(n1705), .B(n1668), .Z(n1242) );
  CENX1 U1833 ( .A(n1704), .B(n1667), .Z(n1243) );
  CENX1 U1834 ( .A(n1621), .B(n1658), .Z(n1180) );
  CENX1 U1835 ( .A(n1622), .B(n1660), .Z(n1178) );
  CENX1 U1836 ( .A(n1622), .B(n1659), .Z(n1179) );
  CENX1 U1837 ( .A(n1698), .B(n1670), .Z(n1288) );
  CENX1 U1838 ( .A(n1704), .B(n1664), .Z(n1246) );
  CENX1 U1839 ( .A(n1705), .B(n1669), .Z(n1241) );
  CENX1 U1840 ( .A(n1658), .B(n1672), .Z(n1167) );
  CENX1 U1841 ( .A(n1617), .B(n1658), .Z(n1300) );
  CENX1 U1842 ( .A(n1617), .B(n1657), .Z(n1301) );
  CENX1 U1843 ( .A(n1709), .B(n1667), .Z(n1222) );
  CENX1 U1844 ( .A(n1621), .B(n1663), .Z(n1175) );
  CENX1 U1845 ( .A(n1658), .B(n1673), .Z(n1156) );
  CENX1 U1846 ( .A(n1659), .B(n1673), .Z(n1155) );
  CENX1 U1847 ( .A(n1567), .B(n1670), .Z(n1408) );
  CENX1 U1848 ( .A(n1657), .B(n1673), .Z(n1157) );
  CENX1 U1849 ( .A(n1660), .B(n1673), .Z(n1154) );
  CENX1 U1850 ( .A(n1661), .B(n1673), .Z(n1153) );
  CENX1 U1851 ( .A(n1678), .B(n1662), .Z(n1416) );
  CENX1 U1852 ( .A(n1567), .B(n1668), .Z(n1410) );
  CENX1 U1853 ( .A(n1567), .B(n1667), .Z(n1411) );
  CENX1 U1854 ( .A(n1687), .B(n1657), .Z(n1357) );
  CENX1 U1855 ( .A(n1709), .B(n1668), .Z(n1221) );
  CENX1 U1856 ( .A(n1682), .B(n1669), .Z(n1376) );
  CENX1 U1857 ( .A(n1704), .B(n1665), .Z(n1245) );
  CENX1 U1858 ( .A(n1705), .B(n1670), .Z(n1240) );
  CENX1 U1859 ( .A(n1672), .B(n1663), .Z(n1162) );
  CENX1 U1860 ( .A(n1680), .B(n1667), .Z(n1378) );
  CENX1 U1861 ( .A(n1662), .B(n1672), .Z(n1163) );
  CENX1 U1862 ( .A(n1704), .B(n1660), .Z(n1250) );
  CENX1 U1863 ( .A(n1704), .B(n1666), .Z(n1244) );
  CENX1 U1864 ( .A(n1702), .B(n1669), .Z(n1264) );
  CENX1 U1865 ( .A(n1680), .B(n1664), .Z(n1381) );
  CENX1 U1866 ( .A(n1674), .B(n1682), .Z(n1390) );
  CENX1 U1867 ( .A(n1674), .B(n1699), .Z(n1303) );
  CENX1 U1868 ( .A(n1674), .B(n1717), .Z(n1198) );
  CENX1 U1869 ( .A(n1674), .B(n1622), .Z(n1183) );
  CENX1 U1870 ( .A(n1661), .B(n1672), .Z(n1164) );
  CENX1 U1871 ( .A(n1682), .B(n1670), .Z(n1375) );
  CENX1 U1872 ( .A(n1716), .B(n1661), .Z(n1192) );
  CENX1 U1873 ( .A(n1716), .B(n1659), .Z(n1194) );
  CENX1 U1874 ( .A(n1660), .B(n1672), .Z(n1165) );
  CENX1 U1875 ( .A(n1709), .B(n1669), .Z(n1220) );
  CENX1 U1876 ( .A(n1713), .B(n1667), .Z(n1203) );
  CENX1 U1877 ( .A(n1713), .B(n1662), .Z(n1208) );
  CENX1 U1878 ( .A(n1682), .B(n1661), .Z(n1384) );
  CENX1 U1879 ( .A(n1565), .B(n1658), .Z(n1356) );
  CENX1 U1880 ( .A(n1680), .B(n1662), .Z(n1383) );
  CENX1 U1881 ( .A(n1683), .B(n1663), .Z(n1382) );
  CENX1 U1882 ( .A(n1674), .B(n1686), .Z(n1359) );
  CIVX2 U1883 ( .A(n1720), .Z(n1717) );
  CENX1 U1884 ( .A(n1675), .B(n1705), .Z(n1255) );
  CNR2IX1 U1885 ( .B(n1675), .A(n114), .Z(n867) );
  CFA1X1 U1886 ( .A(n884), .B(n1028), .CI(n962), .CO(n580), .S(n581) );
  CEOX1 U1887 ( .A(n872), .B(n886), .Z(n429) );
  CENX1 U1888 ( .A(n1680), .B(b[29]), .Z(n1361) );
  CENX1 U1889 ( .A(n1565), .B(b[27]), .Z(n1332) );
  CENX1 U1890 ( .A(n1692), .B(n154), .Z(n1310) );
  CENX1 U1891 ( .A(n1691), .B(n156), .Z(n1308) );
  CENX1 U1892 ( .A(n1691), .B(n157), .Z(n1307) );
  CENX1 U1893 ( .A(n1696), .B(n156), .Z(n1281) );
  CENX1 U1894 ( .A(n1691), .B(b[24]), .Z(n1306) );
  CENX1 U1895 ( .A(n104), .B(a[28]), .Z(n110) );
  CENX1 U1896 ( .A(n1683), .B(n155), .Z(n1369) );
  CENX1 U1897 ( .A(n1698), .B(n157), .Z(n1280) );
  CENX1 U1898 ( .A(n1682), .B(n153), .Z(n1371) );
  CENX1 U1899 ( .A(n1563), .B(b[25]), .Z(n1305) );
  CENX1 U1900 ( .A(n1687), .B(b[25]), .Z(n1334) );
  CENX1 U1901 ( .A(n1686), .B(b[26]), .Z(n1333) );
  CENX1 U1902 ( .A(n1680), .B(n157), .Z(n1367) );
  CENX1 U1903 ( .A(n1657), .B(n104), .Z(n1148) );
  CENX1 U1904 ( .A(n1678), .B(n153), .Z(n1404) );
  CENX1 U1905 ( .A(n1678), .B(n155), .Z(n1402) );
  CENX1 U1906 ( .A(n1678), .B(b[26]), .Z(n1397) );
  CENX1 U1907 ( .A(n1678), .B(b[27]), .Z(n1396) );
  CENX1 U1908 ( .A(n1658), .B(n104), .Z(n1147) );
  CENX1 U1909 ( .A(n1678), .B(n156), .Z(n1401) );
  CENX1 U1910 ( .A(n1678), .B(n157), .Z(n1400) );
  CENX1 U1911 ( .A(n1678), .B(b[25]), .Z(n1398) );
  CENX1 U1912 ( .A(n1678), .B(b[24]), .Z(n1399) );
  CENX1 U1913 ( .A(n1678), .B(b[28]), .Z(n1395) );
  CENX1 U1914 ( .A(n1678), .B(b[29]), .Z(n1394) );
  CENX1 U1915 ( .A(n1678), .B(b[30]), .Z(n1393) );
  CENX1 U1916 ( .A(n1680), .B(n156), .Z(n1368) );
  CENX1 U1917 ( .A(n1660), .B(n104), .Z(n1145) );
  CENX1 U1918 ( .A(n1674), .B(n104), .Z(n1150) );
  CENX1 U1919 ( .A(n1680), .B(b[26]), .Z(n1364) );
  CENX1 U1920 ( .A(n1680), .B(b[27]), .Z(n1363) );
  CENX1 U1921 ( .A(n1684), .B(b[28]), .Z(n1362) );
  CND2X2 U1922 ( .A(n89), .B(n1448), .Z(n91) );
  CND2X1 U1923 ( .A(n1445), .B(n105), .Z(n107) );
  CNIVX2 U1924 ( .A(n116), .Z(n1674) );
  CNIVX4 U1925 ( .A(n99), .Z(n1673) );
  CIVX2 U1926 ( .A(n79), .Z(n1719) );
  CNIVX2 U1927 ( .A(n136), .Z(n1664) );
  CNIVX4 U1928 ( .A(n9), .Z(n1654) );
  CNIVX2 U1929 ( .A(n142), .Z(n1667) );
  CNIVX2 U1930 ( .A(n146), .Z(n1669) );
  CNIVX2 U1931 ( .A(n144), .Z(n1668) );
  CEOX1 U1932 ( .A(a[30]), .B(n113), .Z(n1443) );
  CENX1 U1933 ( .A(n1674), .B(n113), .Z(n1138) );
  CFA1X1 U1935 ( .A(n907), .B(n933), .CI(n919), .CO(n686), .S(n687) );
  CNIVX1 U1936 ( .A(n934), .Z(n1644) );
  COND2XL U1937 ( .A(n97), .B(n1162), .C(n1161), .D(n95), .Z(n886) );
  COND2XL U1938 ( .A(n97), .B(n1164), .C(n1163), .D(n95), .Z(n888) );
  COND2XL U1939 ( .A(n97), .B(n1165), .C(n1164), .D(n95), .Z(n889) );
  COND2XL U1940 ( .A(n97), .B(n1166), .C(n1165), .D(n95), .Z(n890) );
  CNIVX1 U1941 ( .A(n1083), .Z(n1645) );
  CEOX2 U1942 ( .A(a[14]), .B(n1710), .Z(n1451) );
  COND2XL U1943 ( .A(n53), .B(n1258), .C(n1257), .D(n50), .Z(n976) );
  COND2XL U1944 ( .A(n53), .B(n1259), .C(n1258), .D(n50), .Z(n977) );
  COND2XL U1945 ( .A(n53), .B(n1261), .C(n1260), .D(n50), .Z(n979) );
  COND2XL U1946 ( .A(n53), .B(n1265), .C(n1264), .D(n50), .Z(n983) );
  CNR2IX1 U1947 ( .B(n1675), .A(n50), .Z(n997) );
  COND2XL U1948 ( .A(n53), .B(n1276), .C(n1275), .D(n50), .Z(n994) );
  COND2XL U1949 ( .A(n53), .B(n1271), .C(n1270), .D(n50), .Z(n989) );
  CFA1XL U1950 ( .A(n870), .B(n1024), .CI(n958), .CO(n478), .S(n479) );
  COND2X1 U1951 ( .A(n85), .B(n1197), .C(n1196), .D(n82), .Z(n919) );
  COND2XL U1952 ( .A(n77), .B(n1213), .C(n1212), .D(n74), .Z(n934) );
  CIVX1 U1953 ( .A(n1711), .Z(n1710) );
  CIVX2 U1954 ( .A(n1564), .Z(n1689) );
  CIVXL U1955 ( .A(n1564), .Z(n1687) );
  CENX1 U1956 ( .A(n1688), .B(n1667), .Z(n1347) );
  CENX1 U1957 ( .A(n1686), .B(n1666), .Z(n1348) );
  CENX1 U1958 ( .A(n1687), .B(n1668), .Z(n1346) );
  CENX1 U1959 ( .A(n1693), .B(n1658), .Z(n1327) );
  CND2X1 U1960 ( .A(n667), .B(n684), .Z(n1647) );
  CND2X1 U1961 ( .A(n684), .B(n682), .Z(n1649) );
  COND2X1 U1962 ( .A(n27), .B(n1355), .C(n1354), .D(n1559), .Z(n1070) );
  CENX1 U1963 ( .A(n1690), .B(n1661), .Z(n1353) );
  CIVX1 U1964 ( .A(n1685), .Z(n1683) );
  CIVX2 U1965 ( .A(n1685), .Z(n1680) );
  CIVX1 U1966 ( .A(n1685), .Z(n1682) );
  CND2XL U1967 ( .A(n1569), .B(n270), .Z(n175) );
  CND2XL U1968 ( .A(n394), .B(n273), .Z(n176) );
  CIVX1 U1969 ( .A(n272), .Z(n394) );
  COND1XL U1970 ( .A(n358), .B(n360), .C(n359), .Z(n1650) );
  COND2XL U1971 ( .A(n61), .B(n1237), .C(n1236), .D(n58), .Z(n956) );
  COND2XL U1972 ( .A(n61), .B(n1238), .C(n1237), .D(n58), .Z(n957) );
  CNR2IXL U1973 ( .B(n1675), .A(n58), .Z(n975) );
  COND2XL U1974 ( .A(n53), .B(n1703), .C(n1279), .D(n50), .Z(n860) );
  COND2XL U1975 ( .A(n61), .B(n1706), .C(n1256), .D(n58), .Z(n859) );
  COND2XL U1976 ( .A(n61), .B(n1240), .C(n1239), .D(n58), .Z(n959) );
  COND2XL U1977 ( .A(n61), .B(n1245), .C(n1244), .D(n58), .Z(n964) );
  COND2XL U1978 ( .A(n61), .B(n1239), .C(n1238), .D(n58), .Z(n958) );
  COND2XL U1979 ( .A(n61), .B(n1255), .C(n1254), .D(n58), .Z(n974) );
  COND2XL U1980 ( .A(n61), .B(n1251), .C(n1250), .D(n58), .Z(n970) );
  CND2XL U1981 ( .A(n390), .B(n240), .Z(n172) );
  CIVX1 U1982 ( .A(n240), .Z(n238) );
  CIVX1 U1983 ( .A(n239), .Z(n390) );
  CND2XL U1984 ( .A(n391), .B(n250), .Z(n173) );
  CENX1 U1985 ( .A(n1694), .B(n1665), .Z(n1320) );
  CENX1 U1986 ( .A(n1675), .B(n1713), .Z(n1215) );
  CANR1XL U1987 ( .A(n320), .B(n329), .C(n321), .Z(n319) );
  CFA1XL U1988 ( .A(n1015), .B(n1123), .CI(n1065), .CO(n774), .S(n775) );
  CFA1XL U1989 ( .A(n897), .B(n999), .CI(n923), .CO(n452), .S(n453) );
  CNR2X1 U1990 ( .A(n651), .B(n670), .Z(n272) );
  COND2X1 U1991 ( .A(n18), .B(n1370), .C(n1369), .D(n15), .Z(n1084) );
  CENX1 U1992 ( .A(n1680), .B(n154), .Z(n1370) );
  CIVX1 U1993 ( .A(n330), .Z(n329) );
  CENX1 U1994 ( .A(n1690), .B(n156), .Z(n1337) );
  CENX1 U1995 ( .A(n1565), .B(n157), .Z(n1336) );
  COND2XL U1996 ( .A(n69), .B(n1218), .C(n1217), .D(n66), .Z(n938) );
  COND2XL U1997 ( .A(n69), .B(n1219), .C(n1218), .D(n66), .Z(n939) );
  COND2XL U1998 ( .A(n69), .B(n1221), .C(n1220), .D(n66), .Z(n941) );
  COND2XL U1999 ( .A(n69), .B(n1220), .C(n1219), .D(n66), .Z(n940) );
  COND2XL U2000 ( .A(n69), .B(n1711), .C(n1235), .D(n66), .Z(n858) );
  CENX1 U2001 ( .A(n1696), .B(n153), .Z(n1284) );
  CFA1XL U2002 ( .A(n979), .B(n1079), .CI(n1051), .CO(n502), .S(n503) );
  CND2XL U2003 ( .A(n541), .B(n564), .Z(n1651) );
  CND2X1 U2004 ( .A(n541), .B(n543), .Z(n1652) );
  CND2XL U2005 ( .A(n564), .B(n543), .Z(n1653) );
  CND2X1 U2006 ( .A(n513), .B(n538), .Z(n226) );
  CND2X1 U2007 ( .A(n539), .B(n562), .Z(n235) );
  CIVX2 U2008 ( .A(n12), .Z(n1685) );
  CND2IXL U2009 ( .B(n1675), .A(n1683), .Z(n1391) );
  CENXL U2010 ( .A(n1697), .B(n1660), .Z(n1298) );
  CENX1 U2011 ( .A(n1698), .B(n1665), .Z(n1293) );
  CENX1 U2012 ( .A(n1698), .B(n1666), .Z(n1292) );
  CENX1 U2013 ( .A(n1698), .B(n1668), .Z(n1290) );
  CND2IXL U2014 ( .B(n1675), .A(n1690), .Z(n1360) );
  CIVXL U2015 ( .A(n292), .Z(n291) );
  COND1XL U2016 ( .A(n298), .B(n311), .C(n299), .Z(n297) );
  COND2X1 U2017 ( .A(n77), .B(n1214), .C(n1213), .D(n74), .Z(n935) );
  COND2X1 U2018 ( .A(n77), .B(n1206), .C(n1205), .D(n74), .Z(n927) );
  COND2X1 U2019 ( .A(n77), .B(n1207), .C(n1206), .D(n74), .Z(n928) );
  COND2X1 U2020 ( .A(n77), .B(n1205), .C(n1204), .D(n74), .Z(n926) );
  CENX4 U2021 ( .A(n1707), .B(a[16]), .Z(n74) );
  CENX1 U2022 ( .A(n1698), .B(n1667), .Z(n1291) );
  COND2X1 U2023 ( .A(n77), .B(n1210), .C(n1209), .D(n74), .Z(n931) );
  COND2XL U2024 ( .A(n36), .B(n1562), .C(n1331), .D(n1655), .Z(n862) );
  CND2IXL U2025 ( .B(n1675), .A(n1691), .Z(n1331) );
  CENX1 U2026 ( .A(n1691), .B(n153), .Z(n1311) );
  COND2XL U2027 ( .A(n27), .B(n1333), .C(n1332), .D(n1559), .Z(n1048) );
  COND2XL U2028 ( .A(n27), .B(n1352), .C(n1351), .D(n1559), .Z(n1067) );
  COND2XL U2029 ( .A(n27), .B(n1335), .C(n1334), .D(n1559), .Z(n1050) );
  COND2XL U2030 ( .A(n27), .B(n1334), .C(n1333), .D(n1559), .Z(n1049) );
  COND2XL U2031 ( .A(n27), .B(n1359), .C(n1358), .D(n1559), .Z(n1074) );
  COND2XL U2032 ( .A(n27), .B(n1346), .C(n1345), .D(n1559), .Z(n1061) );
  COND2XL U2033 ( .A(n27), .B(n1357), .C(n1356), .D(n1559), .Z(n1072) );
  COND2XL U2034 ( .A(n27), .B(n1354), .C(n1353), .D(n1559), .Z(n1069) );
  COND2XL U2035 ( .A(n27), .B(n1353), .C(n1352), .D(n1559), .Z(n1068) );
  COND2XL U2036 ( .A(n27), .B(n1349), .C(n1348), .D(n1559), .Z(n1064) );
  COND2XL U2037 ( .A(n27), .B(n1356), .C(n1355), .D(n1559), .Z(n1071) );
  COND2XL U2038 ( .A(n27), .B(n1564), .C(n1360), .D(n1559), .Z(n863) );
  COND2XL U2039 ( .A(n27), .B(n1347), .C(n1346), .D(n1559), .Z(n1062) );
  CNR2IXL U2040 ( .B(n1675), .A(n1559), .Z(n1075) );
  COND2XL U2041 ( .A(n27), .B(n1336), .C(n1335), .D(n1559), .Z(n1051) );
  COND2XL U2042 ( .A(n27), .B(n1350), .C(n1349), .D(n1559), .Z(n1065) );
  COND2XL U2043 ( .A(n27), .B(n1358), .C(n1357), .D(n1559), .Z(n1073) );
  COND2XL U2044 ( .A(n27), .B(n1344), .C(n1343), .D(n1559), .Z(n1059) );
  COND2XL U2045 ( .A(n27), .B(n1351), .C(n1350), .D(n1559), .Z(n1066) );
  CENX1 U2046 ( .A(n1698), .B(n1669), .Z(n1289) );
  CIVXL U2047 ( .A(n218), .Z(n387) );
  COND2XL U2048 ( .A(n18), .B(n1362), .C(n1361), .D(n15), .Z(n1076) );
  COND2XL U2049 ( .A(n18), .B(n1363), .C(n1362), .D(n15), .Z(n1077) );
  COND2XL U2050 ( .A(n18), .B(n1364), .C(n1363), .D(n15), .Z(n1078) );
  COND2XL U2051 ( .A(n18), .B(n1388), .C(n1387), .D(n15), .Z(n1102) );
  COND2XL U2052 ( .A(n18), .B(n1386), .C(n1385), .D(n15), .Z(n1100) );
  COND2XL U2053 ( .A(n18), .B(n1385), .C(n1384), .D(n15), .Z(n1099) );
  COND2XL U2054 ( .A(n18), .B(n1383), .C(n1382), .D(n15), .Z(n1097) );
  COND2XL U2055 ( .A(n18), .B(n1382), .C(n1381), .D(n15), .Z(n1096) );
  COND2XL U2056 ( .A(n18), .B(n1366), .C(n1365), .D(n15), .Z(n1080) );
  COND2XL U2057 ( .A(n18), .B(n1379), .C(n1378), .D(n15), .Z(n1093) );
  COND2XL U2058 ( .A(n18), .B(n1384), .C(n1383), .D(n15), .Z(n1098) );
  COND2XL U2059 ( .A(n18), .B(n1365), .C(n1364), .D(n15), .Z(n1079) );
  COND2XL U2060 ( .A(n18), .B(n1369), .C(n1368), .D(n15), .Z(n1083) );
  COND2XL U2061 ( .A(n18), .B(n1685), .C(n1391), .D(n15), .Z(n864) );
  COND2XL U2062 ( .A(n18), .B(n1390), .C(n1389), .D(n15), .Z(n1104) );
  COND2XL U2063 ( .A(n18), .B(n1375), .C(n1374), .D(n15), .Z(n1089) );
  COND2XL U2064 ( .A(n18), .B(n1376), .C(n1375), .D(n15), .Z(n1090) );
  COND2XL U2065 ( .A(n18), .B(n1380), .C(n1379), .D(n15), .Z(n1094) );
  COND2XL U2066 ( .A(n18), .B(n1372), .C(n1371), .D(n15), .Z(n1086) );
  COND2XL U2067 ( .A(n18), .B(n1374), .C(n1373), .D(n15), .Z(n1088) );
  CEOX1 U2068 ( .A(a[2]), .B(n1681), .Z(n1457) );
  CND2X1 U2069 ( .A(n487), .B(n512), .Z(n219) );
  CEOXL U2070 ( .A(n190), .B(n360), .Z(product[7]) );
  CIVX1 U2071 ( .A(n1715), .Z(n1713) );
  COND1XL U2072 ( .A(n261), .B(n278), .C(n262), .Z(n260) );
  CEOXL U2073 ( .A(n236), .B(n171), .Z(product[26]) );
  CENXL U2074 ( .A(n1690), .B(n1665), .Z(n1349) );
  CANR1X2 U2075 ( .A(n312), .B(n293), .C(n294), .Z(n292) );
  COND1X2 U2076 ( .A(n280), .B(n292), .C(n281), .Z(n279) );
  COND2XL U2077 ( .A(n77), .B(n1201), .C(n1200), .D(n74), .Z(n922) );
  COND2XL U2078 ( .A(n77), .B(n1204), .C(n1203), .D(n74), .Z(n925) );
  COND2XL U2079 ( .A(n77), .B(n1203), .C(n1202), .D(n74), .Z(n924) );
  CNR2IXL U2080 ( .B(n1675), .A(n74), .Z(n937) );
  COND2XL U2081 ( .A(n77), .B(n1209), .C(n1208), .D(n74), .Z(n930) );
  COND2XL U2082 ( .A(n77), .B(n1215), .C(n1214), .D(n74), .Z(n936) );
  COND2XL U2083 ( .A(n77), .B(n1202), .C(n1201), .D(n74), .Z(n923) );
  COND2XL U2084 ( .A(n77), .B(n1715), .C(n74), .D(n1216), .Z(n857) );
  CND2IXL U2085 ( .B(n1675), .A(n1707), .Z(n1235) );
  CANR1X2 U2086 ( .A(n275), .B(n1569), .C(n268), .Z(n262) );
  CIVX1 U2087 ( .A(n273), .Z(n275) );
  CEOXL U2088 ( .A(n208), .B(n167), .Z(product[30]) );
  COND2XL U2089 ( .A(n85), .B(n1186), .C(n1185), .D(n82), .Z(n908) );
  COND2XL U2090 ( .A(n85), .B(n1189), .C(n1188), .D(n82), .Z(n911) );
  COND2XL U2091 ( .A(n85), .B(n1188), .C(n1187), .D(n82), .Z(n910) );
  COND2XL U2092 ( .A(n85), .B(n1187), .C(n1186), .D(n82), .Z(n909) );
  COND2XL U2093 ( .A(n85), .B(n1191), .C(n1190), .D(n82), .Z(n913) );
  COND2XL U2094 ( .A(n85), .B(n1190), .C(n1189), .D(n82), .Z(n912) );
  COND2XL U2095 ( .A(n85), .B(n1193), .C(n1192), .D(n82), .Z(n915) );
  COND2XL U2096 ( .A(n85), .B(n1719), .C(n82), .D(n1199), .Z(n856) );
  COND2XL U2097 ( .A(n1198), .B(n85), .C(n1197), .D(n82), .Z(n920) );
  CND2IXL U2098 ( .B(n1675), .A(n1712), .Z(n1216) );
  CENX4 U2099 ( .A(n1679), .B(a[2]), .Z(n15) );
  CND2X4 U2100 ( .A(n1457), .B(n15), .Z(n18) );
  CND2X4 U2101 ( .A(n1453), .B(n50), .Z(n53) );
  CENX4 U2102 ( .A(n1701), .B(a[12]), .Z(n58) );
  CND2X4 U2103 ( .A(n1452), .B(n58), .Z(n61) );
  CENX4 U2104 ( .A(n1704), .B(a[14]), .Z(n66) );
  CND2X4 U2105 ( .A(n1451), .B(n66), .Z(n69) );
  CIVXL U2106 ( .A(n1685), .Z(n1684) );
  CIVXL U2107 ( .A(n1564), .Z(n1686) );
  CIVXL U2108 ( .A(n1564), .Z(n1688) );
  CIVXL U2109 ( .A(n1564), .Z(n1690) );
  CIVXL U2110 ( .A(n1562), .Z(n1692) );
  CIVXL U2111 ( .A(n1562), .Z(n1693) );
  CIVXL U2112 ( .A(n1562), .Z(n1694) );
  CIVXL U2113 ( .A(n1562), .Z(n1695) );
  CIVXL U2114 ( .A(n1700), .Z(n1696) );
  CIVXL U2115 ( .A(n1700), .Z(n1697) );
  CIVXL U2116 ( .A(n1715), .Z(n1714) );
  CIVX2 U2117 ( .A(n374), .Z(n412) );
  CIVX2 U2118 ( .A(n366), .Z(n410) );
  CIVX2 U2119 ( .A(n336), .Z(n404) );
  CIVX2 U2120 ( .A(n333), .Z(n403) );
  CIVX2 U2121 ( .A(n322), .Z(n401) );
  CIVX2 U2122 ( .A(n295), .Z(n397) );
  CIVX2 U2123 ( .A(n234), .Z(n389) );
  CIVX2 U2124 ( .A(n223), .Z(n388) );
  CIVX2 U2125 ( .A(n383), .Z(n381) );
  CIVX2 U2126 ( .A(n380), .Z(n378) );
  CIVX2 U2127 ( .A(n372), .Z(n370) );
  CIVX2 U2128 ( .A(n364), .Z(n362) );
  CIVX2 U2129 ( .A(n356), .Z(n354) );
  CIVX2 U2130 ( .A(n352), .Z(n351) );
  CIVX2 U2131 ( .A(n350), .Z(n348) );
  CIVX2 U2132 ( .A(n345), .Z(n343) );
  CIVX2 U2133 ( .A(n328), .Z(n326) );
  CIVX2 U2134 ( .A(n327), .Z(n402) );
  CIVX2 U2135 ( .A(n312), .Z(n311) );
  CIVX2 U2136 ( .A(n306), .Z(n308) );
  CIVX2 U2137 ( .A(n305), .Z(n399) );
  CIVX2 U2138 ( .A(n303), .Z(n301) );
  CIVX2 U2139 ( .A(n290), .Z(n288) );
  CIVX2 U2140 ( .A(n270), .Z(n268) );
  CIVX2 U2141 ( .A(n261), .Z(n263) );
  CIVX2 U2142 ( .A(n259), .Z(n257) );
  CIVX2 U2143 ( .A(n249), .Z(n391) );
  CIVX2 U2144 ( .A(n212), .Z(n210) );
  CIVX2 U2145 ( .A(n207), .Z(n205) );
  CIVX2 U2146 ( .A(n1621), .Z(n1473) );
  CIVX2 U2147 ( .A(n1672), .Z(n1472) );
  CIVX2 U2148 ( .A(n1673), .Z(n1471) );
  CIVX2 U2149 ( .A(n104), .Z(n1470) );
  CIVX2 U2150 ( .A(n113), .Z(n1468) );
endmodule


module calc_DW_mult_uns_15 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n3, n6, n9, n12, n15, n18, n21, n24, n27, n30, n33, n36, n39, n42,
         n44, n48, n50, n53, n55, n61, n63, n66, n69, n71, n77, n79, n82, n85,
         n87, n89, n91, n93, n95, n97, n99, n100, n102, n104, n105, n107, n109,
         n110, n112, n113, n114, n115, n116, n120, n122, n124, n126, n128,
         n130, n132, n134, n136, n138, n140, n142, n144, n146, n148, n150,
         n151, n152, n153, n154, n155, n156, n157, n166, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n198,
         n199, n205, n206, n207, n208, n210, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n226, n227, n228, n229,
         n231, n234, n235, n236, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n249, n250, n251, n252, n253, n257, n258, n259, n260,
         n261, n262, n263, n264, n268, n270, n271, n272, n273, n275, n278,
         n279, n280, n281, n283, n285, n286, n288, n290, n292, n293, n294,
         n295, n296, n297, n298, n299, n301, n303, n304, n305, n306, n308,
         n311, n312, n313, n314, n316, n318, n319, n320, n321, n322, n323,
         n324, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n343, n345, n346, n348, n350,
         n351, n352, n354, n356, n357, n358, n359, n360, n362, n364, n365,
         n366, n367, n368, n370, n372, n373, n374, n375, n376, n378, n380,
         n381, n383, n385, n387, n388, n389, n390, n391, n392, n394, n397,
         n399, n401, n402, n403, n404, n408, n412, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1451, n1452, n1454, n1455, n1456, n1457, n1458, n1468, n1469, n1470,
         n1471, n1472, n1475, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698;
  assign n3 = a[1];
  assign n12 = a[3];
  assign n21 = a[5];
  assign n30 = a[7];
  assign n39 = a[9];
  assign n48 = a[11];
  assign n55 = a[13];
  assign n63 = a[15];
  assign n71 = a[17];
  assign n79 = a[19];
  assign n87 = a[21];
  assign n93 = a[23];
  assign n99 = a[25];
  assign n104 = a[27];
  assign n109 = a[29];
  assign n113 = a[31];
  assign n116 = b[0];
  assign n120 = b[1];
  assign n122 = b[2];
  assign n124 = b[3];
  assign n126 = b[4];
  assign n128 = b[5];
  assign n130 = b[6];
  assign n132 = b[7];
  assign n134 = b[8];
  assign n136 = b[9];
  assign n138 = b[10];
  assign n140 = b[11];
  assign n142 = b[12];
  assign n144 = b[13];
  assign n146 = b[14];
  assign n148 = b[15];
  assign n150 = b[16];
  assign n151 = b[17];
  assign n152 = b[18];
  assign n153 = b[19];
  assign n154 = b[20];
  assign n155 = b[21];
  assign n156 = b[22];
  assign n157 = b[23];

  CNR2X2 U143 ( .A(n431), .B(n458), .Z(n206) );
  CND2X2 U144 ( .A(n431), .B(n458), .Z(n207) );
  CND2X2 U152 ( .A(n459), .B(n486), .Z(n212) );
  CNR2X2 U183 ( .A(n539), .B(n562), .Z(n234) );
  CEO3X2 U411 ( .A(n422), .B(n421), .C(n440), .Z(n418) );
  CEO3X2 U412 ( .A(n444), .B(n423), .C(n442), .Z(n419) );
  CEO3X2 U413 ( .A(n425), .B(n424), .C(n446), .Z(n420) );
  CEO3X2 U414 ( .A(n428), .B(n427), .C(n426), .Z(n421) );
  CEO3X2 U416 ( .A(n456), .B(n429), .C(n454), .Z(n423) );
  CEO3X2 U417 ( .A(n998), .B(n1106), .C(n1076), .Z(n424) );
  CEO3X2 U418 ( .A(n956), .B(n1048), .C(n866), .Z(n425) );
  CEO3X2 U419 ( .A(n908), .B(n938), .C(n1022), .Z(n426) );
  CEO3X2 U420 ( .A(n896), .B(n922), .C(n976), .Z(n427) );
  CEO3X2 U421 ( .A(n878), .B(n868), .C(n850), .Z(n428) );
  CFA1X1 U423 ( .A(n435), .B(n433), .CI(n460), .CO(n430), .S(n431) );
  CFA1X1 U424 ( .A(n439), .B(n462), .CI(n437), .CO(n432), .S(n433) );
  CFA1X1 U425 ( .A(n441), .B(n464), .CI(n466), .CO(n434), .S(n435) );
  CFA1X1 U426 ( .A(n445), .B(n443), .CI(n468), .CO(n436), .S(n437) );
  CFA1X1 U427 ( .A(n472), .B(n447), .CI(n470), .CO(n438), .S(n439) );
  CFA1X1 U428 ( .A(n451), .B(n449), .CI(n474), .CO(n440), .S(n441) );
  CFA1X1 U429 ( .A(n457), .B(n453), .CI(n455), .CO(n442), .S(n443) );
  CFA1X1 U430 ( .A(n476), .B(n480), .CI(n478), .CO(n444), .S(n445) );
  CFA1X1 U431 ( .A(n1023), .B(n482), .CI(n484), .CO(n446), .S(n447) );
  CFA1X1 U432 ( .A(n957), .B(n1049), .CI(n1107), .CO(n448), .S(n449) );
  CFA1X1 U433 ( .A(n939), .B(n1077), .CI(n999), .CO(n450), .S(n451) );
  CFA1X1 U435 ( .A(n869), .B(n923), .CI(n887), .CO(n454), .S(n455) );
  CFA1X1 U436 ( .A(n867), .B(n879), .CI(n873), .CO(n456), .S(n457) );
  CFA1X1 U437 ( .A(n463), .B(n461), .CI(n488), .CO(n458), .S(n459) );
  CFA1X1 U438 ( .A(n467), .B(n490), .CI(n465), .CO(n460), .S(n461) );
  CFA1X1 U439 ( .A(n469), .B(n492), .CI(n494), .CO(n462), .S(n463) );
  CFA1X1 U440 ( .A(n473), .B(n471), .CI(n496), .CO(n464), .S(n465) );
  CFA1X1 U441 ( .A(n475), .B(n498), .CI(n500), .CO(n466), .S(n467) );
  CFA1X1 U442 ( .A(n481), .B(n477), .CI(n479), .CO(n468), .S(n469) );
  CFA1X1 U443 ( .A(n502), .B(n483), .CI(n504), .CO(n470), .S(n471) );
  CFA1X1 U444 ( .A(n510), .B(n506), .CI(n508), .CO(n472), .S(n473) );
  CFA1X1 U445 ( .A(n1024), .B(n485), .CI(n1108), .CO(n474), .S(n475) );
  CFA1X1 U446 ( .A(n958), .B(n1078), .CI(n1050), .CO(n476), .S(n477) );
  CFA1X1 U449 ( .A(n874), .B(n910), .CI(n898), .CO(n482), .S(n483) );
  CHA1X1 U450 ( .A(n880), .B(n888), .CO(n484), .S(n485) );
  CFA1X1 U451 ( .A(n491), .B(n489), .CI(n514), .CO(n486), .S(n487) );
  CFA1X1 U452 ( .A(n495), .B(n516), .CI(n493), .CO(n488), .S(n489) );
  CFA1X1 U453 ( .A(n497), .B(n518), .CI(n520), .CO(n490), .S(n491) );
  CFA1X1 U454 ( .A(n522), .B(n501), .CI(n499), .CO(n492), .S(n493) );
  CFA1X1 U455 ( .A(n503), .B(n524), .CI(n526), .CO(n494), .S(n495) );
  CFA1X1 U456 ( .A(n509), .B(n505), .CI(n507), .CO(n496), .S(n497) );
  CFA1X1 U457 ( .A(n530), .B(n511), .CI(n528), .CO(n498), .S(n499) );
  CFA1X1 U458 ( .A(n536), .B(n534), .CI(n532), .CO(n500), .S(n501) );
  CFA1X1 U459 ( .A(n979), .B(n1109), .CI(n1001), .CO(n502), .S(n503) );
  CFA1X1 U460 ( .A(n959), .B(n1079), .CI(n1051), .CO(n504), .S(n505) );
  CFA1X1 U461 ( .A(n911), .B(n1025), .CI(n925), .CO(n506), .S(n507) );
  CFA1X1 U462 ( .A(n1589), .B(n941), .CI(n899), .CO(n508), .S(n509) );
  CFA1X1 U463 ( .A(n871), .B(n875), .CI(n881), .CO(n510), .S(n511) );
  CFA1X1 U464 ( .A(n517), .B(n515), .CI(n540), .CO(n512), .S(n513) );
  CFA1X1 U465 ( .A(n521), .B(n542), .CI(n519), .CO(n514), .S(n515) );
  CFA1X1 U466 ( .A(n546), .B(n544), .CI(n523), .CO(n516), .S(n517) );
  CFA1X1 U467 ( .A(n527), .B(n525), .CI(n548), .CO(n518), .S(n519) );
  CFA1X1 U468 ( .A(n535), .B(n550), .CI(n529), .CO(n520), .S(n521) );
  CFA1X1 U469 ( .A(n552), .B(n531), .CI(n533), .CO(n522), .S(n523) );
  CFA1X1 U470 ( .A(n558), .B(n554), .CI(n556), .CO(n524), .S(n525) );
  CFA1X1 U471 ( .A(n1110), .B(n560), .CI(n537), .CO(n526), .S(n527) );
  CFA1X1 U473 ( .A(n942), .B(n876), .CI(n1002), .CO(n530), .S(n531) );
  CFA1X1 U474 ( .A(n852), .B(n960), .CI(n912), .CO(n532), .S(n533) );
  CHA1X1 U476 ( .A(n882), .B(n890), .CO(n536), .S(n537) );
  CFA1X1 U477 ( .A(n543), .B(n541), .CI(n564), .CO(n538), .S(n539) );
  CFA1X1 U478 ( .A(n568), .B(n566), .CI(n545), .CO(n540), .S(n541) );
  CFA1X1 U479 ( .A(n570), .B(n547), .CI(n549), .CO(n542), .S(n543) );
  CFA1X1 U480 ( .A(n574), .B(n551), .CI(n572), .CO(n544), .S(n545) );
  CFA1X1 U481 ( .A(n557), .B(n553), .CI(n555), .CO(n546), .S(n547) );
  CFA1X1 U482 ( .A(n578), .B(n559), .CI(n561), .CO(n548), .S(n549) );
  CFA1X1 U483 ( .A(n582), .B(n576), .CI(n580), .CO(n550), .S(n551) );
  CFA1X1 U484 ( .A(n1003), .B(n584), .CI(n1111), .CO(n552), .S(n553) );
  CFA1X1 U486 ( .A(n1628), .B(n1027), .CI(n943), .CO(n556), .S(n557) );
  CFA1X1 U487 ( .A(n901), .B(n981), .CI(n927), .CO(n558), .S(n559) );
  CFA1X1 U488 ( .A(n877), .B(n891), .CI(n883), .CO(n560), .S(n561) );
  CFA1X1 U489 ( .A(n567), .B(n565), .CI(n588), .CO(n562), .S(n563) );
  CFA1X1 U490 ( .A(n592), .B(n590), .CI(n569), .CO(n564), .S(n565) );
  CFA1X1 U491 ( .A(n594), .B(n571), .CI(n573), .CO(n566), .S(n567) );
  CFA1X1 U492 ( .A(n598), .B(n575), .CI(n596), .CO(n568), .S(n569) );
  CFA1X1 U493 ( .A(n581), .B(n577), .CI(n579), .CO(n570), .S(n571) );
  CFA1X1 U494 ( .A(n602), .B(n583), .CI(n600), .CO(n572), .S(n573) );
  CFA1X1 U495 ( .A(n585), .B(n604), .CI(n606), .CO(n574), .S(n575) );
  CFA1X1 U496 ( .A(n1004), .B(n1082), .CI(n1112), .CO(n576), .S(n577) );
  CFA1X1 U497 ( .A(n962), .B(n884), .CI(n1054), .CO(n578), .S(n579) );
  CFA1X1 U498 ( .A(n914), .B(n1028), .CI(n944), .CO(n580), .S(n581) );
  CFA1X1 U499 ( .A(n902), .B(n928), .CI(n982), .CO(n582), .S(n583) );
  CHA1X1 U500 ( .A(n892), .B(n853), .CO(n584), .S(n585) );
  CFA1X1 U501 ( .A(n591), .B(n589), .CI(n610), .CO(n586), .S(n587) );
  CFA1X1 U502 ( .A(n614), .B(n593), .CI(n612), .CO(n588), .S(n589) );
  CFA1X1 U503 ( .A(n616), .B(n595), .CI(n597), .CO(n590), .S(n591) );
  CFA1X1 U504 ( .A(n620), .B(n599), .CI(n618), .CO(n592), .S(n593) );
  CFA1X1 U505 ( .A(n605), .B(n601), .CI(n603), .CO(n594), .S(n595) );
  CFA1X1 U506 ( .A(n624), .B(n607), .CI(n622), .CO(n596), .S(n597) );
  CFA1X1 U507 ( .A(n1005), .B(n626), .CI(n628), .CO(n598), .S(n599) );
  CFA1X1 U508 ( .A(n983), .B(n1113), .CI(n1055), .CO(n600), .S(n601) );
  CFA1X1 U509 ( .A(n929), .B(n1083), .CI(n963), .CO(n602), .S(n603) );
  CFA1X1 U510 ( .A(n1633), .B(n1029), .CI(n945), .CO(n604), .S(n605) );
  CFA1X1 U511 ( .A(n885), .B(n903), .CI(n893), .CO(n606), .S(n607) );
  CFA1X1 U512 ( .A(n613), .B(n611), .CI(n632), .CO(n608), .S(n609) );
  CFA1X1 U513 ( .A(n617), .B(n634), .CI(n615), .CO(n610), .S(n611) );
  CFA1X1 U515 ( .A(n623), .B(n640), .CI(n621), .CO(n614), .S(n615) );
  CFA1X1 U516 ( .A(n642), .B(n625), .CI(n627), .CO(n616), .S(n617) );
  CFA1X1 U517 ( .A(n648), .B(n644), .CI(n646), .CO(n618), .S(n619) );
  CFA1X1 U518 ( .A(n1114), .B(n629), .CI(n1627), .CO(n620), .S(n621) );
  CFA1X1 U520 ( .A(n916), .B(n1030), .CI(n964), .CO(n624), .S(n625) );
  CFA1X1 U524 ( .A(n639), .B(n654), .CI(n637), .CO(n632), .S(n633) );
  CFA1X1 U525 ( .A(n658), .B(n656), .CI(n641), .CO(n634), .S(n635) );
  CFA1X1 U526 ( .A(n645), .B(n660), .CI(n643), .CO(n636), .S(n637) );
  CFA1X1 U528 ( .A(n668), .B(n664), .CI(n666), .CO(n640), .S(n641) );
  CFA1X1 U529 ( .A(n985), .B(n1115), .CI(n1031), .CO(n642), .S(n643) );
  CFA1X1 U530 ( .A(n947), .B(n1057), .CI(n1007), .CO(n644), .S(n645) );
  CFA1X1 U531 ( .A(n931), .B(n1085), .CI(n965), .CO(n646), .S(n647) );
  CFA1X1 U532 ( .A(n895), .B(n917), .CI(n905), .CO(n648), .S(n649) );
  CFA1X1 U533 ( .A(n655), .B(n653), .CI(n672), .CO(n650), .S(n651) );
  CFA1X1 U534 ( .A(n659), .B(n674), .CI(n657), .CO(n652), .S(n653) );
  CFA1X1 U535 ( .A(n678), .B(n676), .CI(n661), .CO(n654), .S(n655) );
  CFA1X1 U536 ( .A(n665), .B(n663), .CI(n680), .CO(n656), .S(n657) );
  CFA1X1 U537 ( .A(n684), .B(n667), .CI(n682), .CO(n658), .S(n659) );
  CFA1X1 U538 ( .A(n1032), .B(n686), .CI(n669), .CO(n660), .S(n661) );
  CFA1X1 U539 ( .A(n1008), .B(n1116), .CI(n1058), .CO(n662), .S(n663) );
  CFA1X1 U540 ( .A(n855), .B(n1086), .CI(n986), .CO(n664), .S(n665) );
  CFA1X1 U541 ( .A(n932), .B(n906), .CI(n966), .CO(n666), .S(n667) );
  CFA1X1 U543 ( .A(n675), .B(n673), .CI(n690), .CO(n670), .S(n671) );
  CFA1X1 U544 ( .A(n679), .B(n692), .CI(n677), .CO(n672), .S(n673) );
  CFA1X1 U545 ( .A(n681), .B(n694), .CI(n696), .CO(n674), .S(n675) );
  CFA1X1 U546 ( .A(n687), .B(n683), .CI(n685), .CO(n676), .S(n677) );
  CFA1X1 U547 ( .A(n702), .B(n698), .CI(n700), .CO(n678), .S(n679) );
  CFA1X1 U548 ( .A(n987), .B(n704), .CI(n1033), .CO(n680), .S(n681) );
  CFA1X1 U549 ( .A(n967), .B(n1059), .CI(n1117), .CO(n682), .S(n683) );
  CFA1X1 U550 ( .A(n949), .B(n1087), .CI(n1009), .CO(n684), .S(n685) );
  CFA1X1 U551 ( .A(n907), .B(n933), .CI(n919), .CO(n686), .S(n687) );
  CFA1X1 U552 ( .A(n693), .B(n691), .CI(n708), .CO(n688), .S(n689) );
  CFA1X1 U553 ( .A(n697), .B(n710), .CI(n695), .CO(n690), .S(n691) );
  CFA1X1 U554 ( .A(n699), .B(n712), .CI(n714), .CO(n692), .S(n693) );
  CFA1X1 U555 ( .A(n718), .B(n701), .CI(n703), .CO(n694), .S(n695) );
  CFA1X1 U556 ( .A(n705), .B(n716), .CI(n720), .CO(n696), .S(n697) );
  CFA1X1 U557 ( .A(n1034), .B(n1118), .CI(n1060), .CO(n698), .S(n699) );
  CFA1X1 U559 ( .A(n856), .B(n968), .CI(n920), .CO(n702), .S(n703) );
  CHA1X1 U560 ( .A(n934), .B(n988), .CO(n704), .S(n705) );
  CFA1X1 U561 ( .A(n711), .B(n709), .CI(n724), .CO(n706), .S(n707) );
  CFA1X1 U562 ( .A(n715), .B(n726), .CI(n713), .CO(n708), .S(n709) );
  CFA1X1 U563 ( .A(n717), .B(n728), .CI(n730), .CO(n710), .S(n711) );
  CFA1X1 U564 ( .A(n732), .B(n719), .CI(n721), .CO(n712), .S(n713) );
  CFA1X1 U565 ( .A(n1011), .B(n734), .CI(n736), .CO(n714), .S(n715) );
  CFA1X1 U566 ( .A(n989), .B(n1119), .CI(n1035), .CO(n716), .S(n717) );
  CFA1X1 U567 ( .A(n969), .B(n1089), .CI(n1061), .CO(n718), .S(n719) );
  CFA1X1 U568 ( .A(n921), .B(n1637), .CI(n935), .CO(n720), .S(n721) );
  CFA1X1 U569 ( .A(n727), .B(n725), .CI(n740), .CO(n722), .S(n723) );
  CFA1X1 U570 ( .A(n744), .B(n742), .CI(n729), .CO(n724), .S(n725) );
  CFA1X1 U571 ( .A(n735), .B(n731), .CI(n733), .CO(n726), .S(n727) );
  CFA1X1 U572 ( .A(n750), .B(n748), .CI(n746), .CO(n728), .S(n729) );
  CFA1X1 U573 ( .A(n1036), .B(n737), .CI(n1574), .CO(n730), .S(n731) );
  CFA1X1 U574 ( .A(n970), .B(n1090), .CI(n1120), .CO(n732), .S(n733) );
  CFA1X1 U575 ( .A(n952), .B(n936), .CI(n990), .CO(n734), .S(n735) );
  CHA1X1 U576 ( .A(n857), .B(n1012), .CO(n736), .S(n737) );
  CFA1X1 U577 ( .A(n743), .B(n741), .CI(n754), .CO(n738), .S(n739) );
  CFA1X1 U578 ( .A(n758), .B(n756), .CI(n745), .CO(n740), .S(n741) );
  CFA1X1 U579 ( .A(n751), .B(n747), .CI(n749), .CO(n742), .S(n743) );
  CFA1X1 U580 ( .A(n764), .B(n760), .CI(n762), .CO(n744), .S(n745) );
  CFA1X1 U581 ( .A(n1013), .B(n1121), .CI(n1037), .CO(n746), .S(n747) );
  CFA1X1 U582 ( .A(n991), .B(n1091), .CI(n1063), .CO(n748), .S(n749) );
  CFA1X1 U583 ( .A(n937), .B(n971), .CI(n953), .CO(n750), .S(n751) );
  CFA1X1 U584 ( .A(n757), .B(n755), .CI(n768), .CO(n752), .S(n753) );
  CFA1X1 U585 ( .A(n772), .B(n759), .CI(n770), .CO(n754), .S(n755) );
  CFA1X1 U586 ( .A(n774), .B(n761), .CI(n763), .CO(n756), .S(n757) );
  CFA1X1 U587 ( .A(n1038), .B(n776), .CI(n765), .CO(n758), .S(n759) );
  CFA1X1 U588 ( .A(n992), .B(n1092), .CI(n1064), .CO(n760), .S(n761) );
  CFA1X1 U589 ( .A(n972), .B(n954), .CI(n1122), .CO(n762), .S(n763) );
  CHA1X1 U590 ( .A(n858), .B(n1014), .CO(n764), .S(n765) );
  CFA1X1 U591 ( .A(n771), .B(n769), .CI(n780), .CO(n766), .S(n767) );
  CFA1X1 U592 ( .A(n775), .B(n782), .CI(n773), .CO(n768), .S(n769) );
  CFA1X1 U593 ( .A(n784), .B(n777), .CI(n786), .CO(n770), .S(n771) );
  CFA1X1 U594 ( .A(n1039), .B(n788), .CI(n1065), .CO(n772), .S(n773) );
  CFA1X1 U595 ( .A(n1015), .B(n1093), .CI(n1123), .CO(n774), .S(n775) );
  CFA1X1 U596 ( .A(n955), .B(n993), .CI(n973), .CO(n776), .S(n777) );
  CFA1X1 U597 ( .A(n783), .B(n781), .CI(n792), .CO(n778), .S(n779) );
  CFA1X1 U598 ( .A(n787), .B(n794), .CI(n785), .CO(n780), .S(n781) );
  CFA1X1 U599 ( .A(n789), .B(n796), .CI(n798), .CO(n782), .S(n783) );
  CFA1X1 U600 ( .A(n1016), .B(n1040), .CI(n1066), .CO(n784), .S(n785) );
  CFA1X1 U601 ( .A(n994), .B(n974), .CI(n1124), .CO(n786), .S(n787) );
  CFA1X1 U603 ( .A(n802), .B(n793), .CI(n795), .CO(n790), .S(n791) );
  CFA1X1 U604 ( .A(n799), .B(n804), .CI(n797), .CO(n792), .S(n793) );
  CFA1X1 U605 ( .A(n1125), .B(n806), .CI(n808), .CO(n794), .S(n795) );
  CFA1X1 U606 ( .A(n1041), .B(n1095), .CI(n1067), .CO(n796), .S(n797) );
  CFA1X1 U607 ( .A(n975), .B(n1017), .CI(n995), .CO(n798), .S(n799) );
  CFA1X1 U608 ( .A(n805), .B(n803), .CI(n812), .CO(n800), .S(n801) );
  CFA1X1 U609 ( .A(n816), .B(n807), .CI(n814), .CO(n802), .S(n803) );
  CFA1X1 U610 ( .A(n1042), .B(n809), .CI(n1068), .CO(n804), .S(n805) );
  CFA1X1 U611 ( .A(n1018), .B(n1096), .CI(n1126), .CO(n806), .S(n807) );
  CHA1X1 U612 ( .A(n860), .B(n996), .CO(n808), .S(n809) );
  CFA1X1 U613 ( .A(n815), .B(n813), .CI(n820), .CO(n810), .S(n811) );
  CFA1X1 U614 ( .A(n824), .B(n817), .CI(n822), .CO(n812), .S(n813) );
  CFA1X1 U615 ( .A(n1127), .B(n1097), .CI(n1069), .CO(n814), .S(n815) );
  CFA1X1 U616 ( .A(n997), .B(n1043), .CI(n1019), .CO(n816), .S(n817) );
  CFA1X1 U617 ( .A(n828), .B(n821), .CI(n823), .CO(n818), .S(n819) );
  CFA1X1 U618 ( .A(n1128), .B(n830), .CI(n825), .CO(n820), .S(n821) );
  CFA1X1 U619 ( .A(n1044), .B(n1098), .CI(n1070), .CO(n822), .S(n823) );
  CHA1X1 U620 ( .A(n861), .B(n1020), .CO(n824), .S(n825) );
  CFA1X1 U621 ( .A(n834), .B(n829), .CI(n831), .CO(n826), .S(n827) );
  CFA1X1 U622 ( .A(n1071), .B(n836), .CI(n1099), .CO(n828), .S(n829) );
  CFA1X1 U623 ( .A(n1021), .B(n1129), .CI(n1045), .CO(n830), .S(n831) );
  CFA1X1 U624 ( .A(n837), .B(n835), .CI(n840), .CO(n832), .S(n833) );
  CFA1X1 U625 ( .A(n1130), .B(n1100), .CI(n1072), .CO(n834), .S(n835) );
  CHA1X1 U626 ( .A(n862), .B(n1046), .CO(n836), .S(n837) );
  CFA1X1 U627 ( .A(n1101), .B(n841), .CI(n844), .CO(n838), .S(n839) );
  CFA1X1 U628 ( .A(n1047), .B(n1073), .CI(n1131), .CO(n840), .S(n841) );
  CFA1X1 U629 ( .A(n1132), .B(n845), .CI(n1102), .CO(n842), .S(n843) );
  CHA1X1 U630 ( .A(n863), .B(n1074), .CO(n844), .S(n845) );
  CHA1X1 U632 ( .A(n1134), .B(n864), .CO(n848), .S(n849) );
  COND2X1 U633 ( .A(n1139), .B(n114), .C(n1468), .D(n115), .Z(n850) );
  COND2X1 U634 ( .A(n1138), .B(n115), .C(n114), .D(n1137), .Z(n866) );
  CND2IX1 U638 ( .B(n1559), .A(n113), .Z(n1139) );
  COND2X1 U639 ( .A(n1144), .B(n110), .C(n1469), .D(n112), .Z(n851) );
  COND2X1 U640 ( .A(n112), .B(n1141), .C(n110), .D(n1140), .Z(n868) );
  COND2X1 U641 ( .A(n112), .B(n1142), .C(n110), .D(n1141), .Z(n869) );
  COND2X1 U642 ( .A(n1143), .B(n112), .C(n110), .D(n1142), .Z(n870) );
  COND2X1 U650 ( .A(n107), .B(n1146), .C(n105), .D(n1145), .Z(n872) );
  COND2X1 U651 ( .A(n107), .B(n1147), .C(n105), .D(n1146), .Z(n873) );
  COND2X1 U652 ( .A(n107), .B(n1148), .C(n105), .D(n1147), .Z(n874) );
  COND2X1 U653 ( .A(n1149), .B(n107), .C(n105), .D(n1148), .Z(n875) );
  COND2X1 U654 ( .A(n1150), .B(n107), .C(n105), .D(n1149), .Z(n876) );
  CND2IX1 U662 ( .B(n1559), .A(n104), .Z(n1151) );
  COND2X1 U663 ( .A(n1160), .B(n1592), .C(n1471), .D(n102), .Z(n853) );
  COND2X1 U664 ( .A(n102), .B(n1153), .C(n1592), .D(n1152), .Z(n878) );
  COND2X1 U665 ( .A(n102), .B(n1154), .C(n1592), .D(n1153), .Z(n879) );
  COND2X1 U666 ( .A(n102), .B(n1155), .C(n1592), .D(n1154), .Z(n880) );
  COND2X1 U667 ( .A(n102), .B(n1156), .C(n1592), .D(n1155), .Z(n881) );
  COND2X1 U668 ( .A(n102), .B(n1157), .C(n1592), .D(n1156), .Z(n882) );
  COND2X1 U669 ( .A(n102), .B(n1158), .C(n1592), .D(n1157), .Z(n883) );
  COND2X1 U670 ( .A(n1159), .B(n102), .C(n1592), .D(n1158), .Z(n884) );
  CND2IX1 U680 ( .B(n1559), .A(n1648), .Z(n1160) );
  COND2X1 U683 ( .A(n97), .B(n1163), .C(n1162), .D(n95), .Z(n887) );
  COND2X1 U687 ( .A(n97), .B(n1167), .C(n95), .D(n1166), .Z(n891) );
  COND2X1 U688 ( .A(n97), .B(n1168), .C(n95), .D(n1167), .Z(n892) );
  COND2X1 U689 ( .A(n97), .B(n1169), .C(n95), .D(n1168), .Z(n893) );
  CND2IX1 U702 ( .B(n1559), .A(n1647), .Z(n1171) );
  COND2X1 U703 ( .A(n1184), .B(n89), .C(n1585), .D(n91), .Z(n855) );
  COND2X1 U709 ( .A(n91), .B(n1178), .C(n1177), .D(n89), .Z(n901) );
  COND2X1 U710 ( .A(n91), .B(n1179), .C(n1178), .D(n89), .Z(n902) );
  COND2X1 U713 ( .A(n91), .B(n1182), .C(n89), .D(n1181), .Z(n905) );
  CND2IX1 U728 ( .B(n1559), .A(n1646), .Z(n1184) );
  COND2X1 U729 ( .A(n85), .B(n1593), .C(n82), .D(n1199), .Z(n856) );
  COND2X1 U734 ( .A(n85), .B(n1190), .C(n1189), .D(n82), .Z(n912) );
  COND2X1 U736 ( .A(n85), .B(n1192), .C(n1191), .D(n82), .Z(n914) );
  COND2X1 U739 ( .A(n85), .B(n1195), .C(n1194), .D(n82), .Z(n917) );
  COND2X1 U740 ( .A(n85), .B(n1196), .C(n1195), .D(n82), .Z(n918) );
  COND2X1 U741 ( .A(n85), .B(n1197), .C(n1196), .D(n82), .Z(n919) );
  COND2X1 U759 ( .A(n77), .B(n1475), .C(n1635), .D(n1216), .Z(n857) );
  COND2X1 U764 ( .A(n77), .B(n1205), .C(n1204), .D(n1635), .Z(n926) );
  COND2X1 U765 ( .A(n77), .B(n1206), .C(n1205), .D(n1635), .Z(n927) );
  COND2X1 U766 ( .A(n77), .B(n1207), .C(n1206), .D(n1635), .Z(n928) );
  COND2X1 U767 ( .A(n77), .B(n1208), .C(n1207), .D(n1635), .Z(n929) );
  COND2X1 U770 ( .A(n77), .B(n1211), .C(n1210), .D(n1635), .Z(n932) );
  COND2X1 U771 ( .A(n77), .B(n1212), .C(n1211), .D(n1635), .Z(n933) );
  COND2X1 U773 ( .A(n77), .B(n1214), .C(n1213), .D(n1635), .Z(n935) );
  COND2X1 U798 ( .A(n69), .B(n1222), .C(n1221), .D(n66), .Z(n942) );
  COND2X1 U800 ( .A(n69), .B(n1224), .C(n1223), .D(n66), .Z(n944) );
  COND2X1 U805 ( .A(n69), .B(n1229), .C(n1228), .D(n66), .Z(n949) );
  COND2X1 U809 ( .A(n69), .B(n1233), .C(n1232), .D(n66), .Z(n953) );
  CND2IX1 U830 ( .B(n1559), .A(n1693), .Z(n1235) );
  COND2X1 U832 ( .A(n61), .B(n1237), .C(n1236), .D(n1630), .Z(n956) );
  COND2X1 U834 ( .A(n61), .B(n1239), .C(n1238), .D(n1631), .Z(n958) );
  COND2X1 U835 ( .A(n61), .B(n1240), .C(n1239), .D(n1630), .Z(n959) );
  COND2X1 U836 ( .A(n61), .B(n1241), .C(n1240), .D(n1631), .Z(n960) );
  COND2X1 U837 ( .A(n61), .B(n1242), .C(n1241), .D(n1631), .Z(n961) );
  COND2X1 U838 ( .A(n61), .B(n1243), .C(n1242), .D(n1631), .Z(n962) );
  COND2X1 U839 ( .A(n61), .B(n1244), .C(n1243), .D(n1630), .Z(n963) );
  COND2X1 U840 ( .A(n61), .B(n1245), .C(n1244), .D(n1630), .Z(n964) );
  COND2X1 U841 ( .A(n61), .B(n1246), .C(n1245), .D(n1631), .Z(n965) );
  COND2X1 U842 ( .A(n61), .B(n1247), .C(n1246), .D(n1631), .Z(n966) );
  COND2X1 U843 ( .A(n61), .B(n1248), .C(n1247), .D(n1630), .Z(n967) );
  COND2X1 U844 ( .A(n61), .B(n1249), .C(n1248), .D(n1630), .Z(n968) );
  COND2X1 U845 ( .A(n61), .B(n1250), .C(n1249), .D(n1631), .Z(n969) );
  COND2X1 U846 ( .A(n61), .B(n1251), .C(n1250), .D(n1630), .Z(n970) );
  COND2X1 U847 ( .A(n61), .B(n1252), .C(n1251), .D(n1631), .Z(n971) );
  COND2X1 U848 ( .A(n61), .B(n1253), .C(n1252), .D(n1631), .Z(n972) );
  COND2X1 U849 ( .A(n61), .B(n1254), .C(n1253), .D(n1631), .Z(n973) );
  COND2X1 U850 ( .A(n1255), .B(n61), .C(n1254), .D(n1630), .Z(n974) );
  COND2X1 U880 ( .A(n53), .B(n1264), .C(n1263), .D(n1597), .Z(n982) );
  COND2X1 U881 ( .A(n53), .B(n1265), .C(n1264), .D(n1597), .Z(n983) );
  COND2X1 U883 ( .A(n53), .B(n1267), .C(n1266), .D(n1597), .Z(n985) );
  COND2X1 U884 ( .A(n53), .B(n1268), .C(n1267), .D(n1597), .Z(n986) );
  COND2X1 U889 ( .A(n53), .B(n1273), .C(n1272), .D(n1597), .Z(n991) );
  COND2X1 U890 ( .A(n53), .B(n1274), .C(n1273), .D(n1597), .Z(n992) );
  COND2X1 U891 ( .A(n53), .B(n1275), .C(n1274), .D(n1597), .Z(n993) );
  COND2X1 U922 ( .A(n44), .B(n1283), .C(n1282), .D(n42), .Z(n1000) );
  COND2X1 U923 ( .A(n44), .B(n1284), .C(n1283), .D(n42), .Z(n1001) );
  COND2X1 U924 ( .A(n44), .B(n1285), .C(n1284), .D(n42), .Z(n1002) );
  COND2X1 U925 ( .A(n44), .B(n1286), .C(n1285), .D(n42), .Z(n1003) );
  COND2X1 U928 ( .A(n44), .B(n1289), .C(n1288), .D(n42), .Z(n1006) );
  COND2X1 U929 ( .A(n44), .B(n1290), .C(n1289), .D(n42), .Z(n1007) );
  COND2X1 U930 ( .A(n44), .B(n1291), .C(n1290), .D(n42), .Z(n1008) );
  COND2X1 U931 ( .A(n44), .B(n1292), .C(n1291), .D(n42), .Z(n1009) );
  COND2X1 U932 ( .A(n44), .B(n1293), .C(n1292), .D(n42), .Z(n1010) );
  COND2X1 U934 ( .A(n44), .B(n1295), .C(n1294), .D(n42), .Z(n1012) );
  COND2X1 U935 ( .A(n44), .B(n1296), .C(n1295), .D(n42), .Z(n1013) );
  COND2X1 U937 ( .A(n44), .B(n1298), .C(n1297), .D(n42), .Z(n1015) );
  COND2X1 U938 ( .A(n44), .B(n1299), .C(n1298), .D(n42), .Z(n1016) );
  COND2X1 U939 ( .A(n44), .B(n1300), .C(n1299), .D(n42), .Z(n1017) );
  COND2X1 U940 ( .A(n44), .B(n1301), .C(n1300), .D(n42), .Z(n1018) );
  COND2X1 U941 ( .A(n44), .B(n1302), .C(n1301), .D(n42), .Z(n1019) );
  COND2X1 U974 ( .A(n36), .B(n1310), .C(n1309), .D(n33), .Z(n1026) );
  COND2X1 U975 ( .A(n36), .B(n1311), .C(n1310), .D(n33), .Z(n1027) );
  COND2X1 U976 ( .A(n36), .B(n1312), .C(n1311), .D(n33), .Z(n1028) );
  COND2X1 U979 ( .A(n36), .B(n1315), .C(n1314), .D(n33), .Z(n1031) );
  COND2X1 U981 ( .A(n36), .B(n1317), .C(n1316), .D(n33), .Z(n1033) );
  COND2X1 U983 ( .A(n36), .B(n1319), .C(n1318), .D(n33), .Z(n1035) );
  COND2X1 U984 ( .A(n36), .B(n1320), .C(n1319), .D(n33), .Z(n1036) );
  COND2X1 U985 ( .A(n36), .B(n1321), .C(n1320), .D(n33), .Z(n1037) );
  COND2X1 U991 ( .A(n36), .B(n1327), .C(n1326), .D(n33), .Z(n1043) );
  COND2X1 U992 ( .A(n36), .B(n1328), .C(n1327), .D(n33), .Z(n1044) );
  COND2X1 U1026 ( .A(n27), .B(n1335), .C(n1334), .D(n24), .Z(n1050) );
  COND2X1 U1028 ( .A(n27), .B(n1337), .C(n1336), .D(n24), .Z(n1052) );
  COND2X1 U1029 ( .A(n27), .B(n1338), .C(n1337), .D(n24), .Z(n1053) );
  COND2X1 U1030 ( .A(n27), .B(n1339), .C(n1338), .D(n24), .Z(n1054) );
  COND2X1 U1031 ( .A(n27), .B(n1340), .C(n1339), .D(n24), .Z(n1055) );
  COND2X1 U1033 ( .A(n27), .B(n1342), .C(n1341), .D(n24), .Z(n1057) );
  COND2X1 U1034 ( .A(n27), .B(n1343), .C(n1342), .D(n24), .Z(n1058) );
  COND2X1 U1035 ( .A(n27), .B(n1344), .C(n1343), .D(n24), .Z(n1059) );
  COND2X1 U1037 ( .A(n27), .B(n1346), .C(n1345), .D(n24), .Z(n1061) );
  COND2X1 U1039 ( .A(n27), .B(n1348), .C(n1347), .D(n24), .Z(n1063) );
  COND2X1 U1040 ( .A(n27), .B(n1349), .C(n1348), .D(n24), .Z(n1064) );
  COND2X1 U1042 ( .A(n27), .B(n1351), .C(n1350), .D(n24), .Z(n1066) );
  COND2X1 U1043 ( .A(n27), .B(n1352), .C(n1351), .D(n24), .Z(n1067) );
  CND2IX1 U1080 ( .B(n1559), .A(n1666), .Z(n1360) );
  COND2X1 U1086 ( .A(n18), .B(n1366), .C(n15), .D(n1365), .Z(n1080) );
  COND2X1 U1088 ( .A(n18), .B(n1368), .C(n15), .D(n1367), .Z(n1082) );
  COND2X1 U1091 ( .A(n18), .B(n1371), .C(n15), .D(n1370), .Z(n1085) );
  COND2X1 U1092 ( .A(n18), .B(n1372), .C(n15), .D(n1371), .Z(n1086) );
  COND2X1 U1093 ( .A(n18), .B(n1373), .C(n15), .D(n1372), .Z(n1087) );
  COND2X1 U1094 ( .A(n18), .B(n1374), .C(n15), .D(n1373), .Z(n1088) );
  COND2X1 U1095 ( .A(n18), .B(n1375), .C(n15), .D(n1374), .Z(n1089) );
  COND2X1 U1097 ( .A(n18), .B(n1377), .C(n15), .D(n1376), .Z(n1091) );
  COND2X1 U1098 ( .A(n18), .B(n1378), .C(n15), .D(n1377), .Z(n1092) );
  COND2X1 U1144 ( .A(n9), .B(n1393), .C(n6), .D(n1392), .Z(n1106) );
  COND2X1 U1145 ( .A(n9), .B(n1394), .C(n6), .D(n1393), .Z(n1107) );
  COND2X1 U1146 ( .A(n9), .B(n1395), .C(n6), .D(n1394), .Z(n1108) );
  COND2X1 U1147 ( .A(n9), .B(n1396), .C(n6), .D(n1395), .Z(n1109) );
  COND2X1 U1148 ( .A(n9), .B(n1397), .C(n6), .D(n1396), .Z(n1110) );
  COND2X1 U1149 ( .A(n9), .B(n1398), .C(n6), .D(n1397), .Z(n1111) );
  COND2X1 U1151 ( .A(n9), .B(n1400), .C(n6), .D(n1399), .Z(n1113) );
  COND2X1 U1152 ( .A(n9), .B(n1401), .C(n6), .D(n1400), .Z(n1114) );
  COND2X1 U1153 ( .A(n9), .B(n1402), .C(n6), .D(n1401), .Z(n1115) );
  COND2X1 U1154 ( .A(n9), .B(n1403), .C(n6), .D(n1402), .Z(n1116) );
  COND2X1 U1155 ( .A(n9), .B(n1404), .C(n6), .D(n1403), .Z(n1117) );
  COND2X1 U1156 ( .A(n9), .B(n1405), .C(n6), .D(n1404), .Z(n1118) );
  COND2X1 U1157 ( .A(n9), .B(n1406), .C(n6), .D(n1405), .Z(n1119) );
  COND2X1 U1158 ( .A(n9), .B(n1407), .C(n6), .D(n1406), .Z(n1120) );
  COND2X1 U1159 ( .A(n9), .B(n1408), .C(n6), .D(n1407), .Z(n1121) );
  COND2X1 U1160 ( .A(n9), .B(n1409), .C(n6), .D(n1408), .Z(n1122) );
  COND2X1 U1161 ( .A(n9), .B(n1410), .C(n6), .D(n1409), .Z(n1123) );
  COND2X1 U1162 ( .A(n9), .B(n1411), .C(n6), .D(n1410), .Z(n1124) );
  COND2X1 U1163 ( .A(n9), .B(n1412), .C(n6), .D(n1411), .Z(n1125) );
  COND2X1 U1164 ( .A(n9), .B(n1413), .C(n6), .D(n1412), .Z(n1126) );
  COND2X1 U1165 ( .A(n9), .B(n1414), .C(n6), .D(n1413), .Z(n1127) );
  COND2X1 U1166 ( .A(n9), .B(n1415), .C(n6), .D(n1414), .Z(n1128) );
  COND2X1 U1167 ( .A(n9), .B(n1416), .C(n6), .D(n1415), .Z(n1129) );
  COND2X1 U1168 ( .A(n9), .B(n1417), .C(n6), .D(n1416), .Z(n1130) );
  COND2X1 U1169 ( .A(n9), .B(n1418), .C(n6), .D(n1417), .Z(n1131) );
  COND2X1 U1170 ( .A(n9), .B(n1419), .C(n6), .D(n1418), .Z(n1132) );
  COND2X1 U1171 ( .A(n9), .B(n1420), .C(n6), .D(n1419), .Z(n1133) );
  COND2X1 U1172 ( .A(n9), .B(n1421), .C(n6), .D(n1420), .Z(n1134) );
  COND2X1 U1173 ( .A(n9), .B(n1422), .C(n6), .D(n1421), .Z(n1135) );
  COND2X1 U1174 ( .A(n1423), .B(n9), .C(n6), .D(n1422), .Z(n1136) );
  CND2X2 U1237 ( .A(n1445), .B(n105), .Z(n107) );
  CEOX2 U1256 ( .A(a[14]), .B(n1697), .Z(n1451) );
  CEOX2 U1259 ( .A(a[12]), .B(n1691), .Z(n1452) );
  CEOX2 U1265 ( .A(a[8]), .B(n1682), .Z(n1454) );
  CEOX2 U1271 ( .A(a[4]), .B(n1672), .Z(n1456) );
  CEOX2 U1274 ( .A(a[2]), .B(n1664), .Z(n1457) );
  COND1XL U1281 ( .A(n214), .B(n242), .C(n1575), .Z(n1557) );
  COND1XL U1282 ( .A(n214), .B(n242), .C(n1575), .Z(n1577) );
  COND1X1 U1283 ( .A(n368), .B(n366), .C(n367), .Z(n365) );
  CND2X4 U1284 ( .A(n89), .B(n1448), .Z(n91) );
  CENXL U1285 ( .A(n1696), .B(n150), .Z(n1218) );
  COND2XL U1286 ( .A(n27), .B(n1345), .C(n1344), .D(n24), .Z(n1060) );
  CNR2X2 U1287 ( .A(n513), .B(n538), .Z(n223) );
  COND2XL U1288 ( .A(n44), .B(n1281), .C(n1280), .D(n42), .Z(n998) );
  COND2XL U1289 ( .A(n44), .B(n1282), .C(n1281), .D(n42), .Z(n999) );
  COND2XL U1290 ( .A(n44), .B(n1294), .C(n1293), .D(n42), .Z(n1011) );
  COND2XL U1291 ( .A(n1303), .B(n44), .C(n1302), .D(n42), .Z(n1020) );
  COND2XL U1292 ( .A(n44), .B(n1288), .C(n1287), .D(n42), .Z(n1005) );
  CENXL U1293 ( .A(n1644), .B(n148), .Z(n1200) );
  CENXL U1294 ( .A(n1559), .B(n1644), .Z(n1215) );
  CENXL U1295 ( .A(n1651), .B(n1644), .Z(n1214) );
  CENXL U1296 ( .A(n1644), .B(n1562), .Z(n1213) );
  CENXL U1297 ( .A(n1644), .B(n142), .Z(n1203) );
  CENXL U1298 ( .A(n1644), .B(n1564), .Z(n1210) );
  CENX1 U1299 ( .A(n1644), .B(n138), .Z(n1205) );
  CFA1XL U1300 ( .A(n1075), .B(n1103), .CI(n1133), .CO(n846), .S(n847) );
  CENXL U1301 ( .A(n1657), .B(b[28]), .Z(n1362) );
  CENX1 U1302 ( .A(n1657), .B(n153), .Z(n1371) );
  CENX1 U1303 ( .A(n1694), .B(n134), .Z(n1226) );
  CENXL U1304 ( .A(n1654), .B(n138), .Z(n1413) );
  CENXL U1305 ( .A(n1645), .B(n138), .Z(n1188) );
  CIVX4 U1306 ( .A(n1698), .Z(n1693) );
  CIVX4 U1307 ( .A(n63), .Z(n1698) );
  CIVX2 U1308 ( .A(n1625), .Z(n1635) );
  CENXL U1309 ( .A(n136), .B(n1647), .Z(n1161) );
  CENXL U1310 ( .A(n1654), .B(n136), .Z(n1414) );
  CENXL U1311 ( .A(n1662), .B(n136), .Z(n1381) );
  CENXL U1312 ( .A(n1644), .B(n136), .Z(n1206) );
  CENXL U1313 ( .A(n1645), .B(n136), .Z(n1189) );
  CNIVXL U1314 ( .A(n1650), .Z(n1558) );
  CNIVX4 U1315 ( .A(n1650), .Z(n1559) );
  CNIVXL U1316 ( .A(n116), .Z(n1650) );
  CENXL U1317 ( .A(n1691), .B(n153), .Z(n1236) );
  CENXL U1318 ( .A(n1653), .B(n153), .Z(n1404) );
  CENXL U1319 ( .A(n132), .B(n1648), .Z(n1152) );
  CENXL U1320 ( .A(n1659), .B(n132), .Z(n1383) );
  CENXL U1321 ( .A(n1668), .B(n132), .Z(n1352) );
  CENXL U1322 ( .A(n1674), .B(n132), .Z(n1323) );
  CENXL U1323 ( .A(n132), .B(n1647), .Z(n1163) );
  CENXL U1324 ( .A(n1681), .B(n132), .Z(n1296) );
  CENXL U1325 ( .A(n1690), .B(n132), .Z(n1248) );
  CENXL U1326 ( .A(n1644), .B(n132), .Z(n1208) );
  CENXL U1327 ( .A(n1645), .B(n132), .Z(n1191) );
  CENXL U1328 ( .A(n1668), .B(n130), .Z(n1353) );
  CENXL U1329 ( .A(n1681), .B(n130), .Z(n1297) );
  CENXL U1330 ( .A(n1654), .B(n130), .Z(n1417) );
  CENXL U1331 ( .A(n1674), .B(n130), .Z(n1324) );
  CENXL U1332 ( .A(n1687), .B(n130), .Z(n1272) );
  CENXL U1333 ( .A(n130), .B(n1648), .Z(n1153) );
  CENXL U1334 ( .A(n1646), .B(n130), .Z(n1177) );
  CENXL U1335 ( .A(n1693), .B(n130), .Z(n1228) );
  CENXL U1336 ( .A(n1644), .B(n130), .Z(n1209) );
  CENXL U1337 ( .A(n1645), .B(n130), .Z(n1192) );
  CENXL U1338 ( .A(n1654), .B(n134), .Z(n1415) );
  CENXL U1339 ( .A(n1662), .B(n134), .Z(n1382) );
  CENXL U1340 ( .A(n1646), .B(n134), .Z(n1175) );
  CENXL U1341 ( .A(n1670), .B(n134), .Z(n1351) );
  CENXL U1342 ( .A(n1674), .B(n134), .Z(n1322) );
  CENXL U1343 ( .A(n1684), .B(n134), .Z(n1295) );
  CENXL U1344 ( .A(n1644), .B(n134), .Z(n1207) );
  CENXL U1345 ( .A(n1646), .B(n140), .Z(n1172) );
  CENXL U1346 ( .A(n1654), .B(n140), .Z(n1412) );
  CENXL U1347 ( .A(n1661), .B(n140), .Z(n1379) );
  CENXL U1348 ( .A(n1670), .B(n140), .Z(n1348) );
  CENXL U1349 ( .A(n1676), .B(n140), .Z(n1319) );
  CENXL U1350 ( .A(n1688), .B(n140), .Z(n1267) );
  CENXL U1351 ( .A(n1645), .B(n140), .Z(n1187) );
  CENXL U1352 ( .A(n1683), .B(n140), .Z(n1292) );
  CIVX3 U1353 ( .A(n55), .Z(n1692) );
  COND2X1 U1354 ( .A(n1151), .B(n105), .C(n1470), .D(n107), .Z(n852) );
  CIVX3 U1355 ( .A(n1665), .Z(n1661) );
  CENX1 U1356 ( .A(n1691), .B(n152), .Z(n1237) );
  CND3X1 U1357 ( .A(n1578), .B(n1579), .C(n1580), .Z(n638) );
  CENX1 U1358 ( .A(n1644), .B(n1563), .Z(n1211) );
  CENX1 U1359 ( .A(n1649), .B(n1645), .Z(n1198) );
  CENX1 U1360 ( .A(n1644), .B(n1561), .Z(n1212) );
  CENX1 U1361 ( .A(n1683), .B(n152), .Z(n1285) );
  CENX1 U1362 ( .A(n1653), .B(b[26]), .Z(n1397) );
  CENX1 U1363 ( .A(n1559), .B(n1691), .Z(n1255) );
  CENX1 U1364 ( .A(n1682), .B(n1561), .Z(n1300) );
  CENX1 U1365 ( .A(n1645), .B(n1564), .Z(n1193) );
  CENX1 U1366 ( .A(n1691), .B(n150), .Z(n1239) );
  CFA1X1 U1367 ( .A(n1052), .B(n1080), .CI(n1026), .CO(n528), .S(n529) );
  CENX1 U1368 ( .A(n1668), .B(n1564), .Z(n1354) );
  CENX1 U1369 ( .A(n1561), .B(n1645), .Z(n1195) );
  CENX1 U1370 ( .A(n1645), .B(n1563), .Z(n1194) );
  CNIVX1 U1371 ( .A(n1084), .Z(n1632) );
  CENX1 U1372 ( .A(n1651), .B(n109), .Z(n1142) );
  CENX1 U1373 ( .A(n1562), .B(n109), .Z(n1141) );
  CIVX2 U1374 ( .A(n1639), .Z(n33) );
  CND2X2 U1375 ( .A(n1454), .B(n42), .Z(n44) );
  CIVX4 U1376 ( .A(n1626), .Z(n42) );
  CEOX2 U1377 ( .A(n30), .B(a[8]), .Z(n1626) );
  CENX1 U1378 ( .A(n1691), .B(n151), .Z(n1238) );
  CND3X1 U1379 ( .A(n1582), .B(n1583), .C(n1584), .Z(n612) );
  CENX1 U1380 ( .A(n1649), .B(n113), .Z(n1138) );
  CEOX1 U1381 ( .A(a[26]), .B(n104), .Z(n1445) );
  CIVX3 U1382 ( .A(n3), .Z(n1656) );
  CENX1 U1383 ( .A(n1649), .B(n1664), .Z(n1390) );
  CANR1XL U1384 ( .A(n348), .B(n1614), .C(n343), .Z(n341) );
  CEOX1 U1385 ( .A(n1581), .B(n638), .Z(n613) );
  COND1X1 U1386 ( .A(n280), .B(n292), .C(n281), .Z(n279) );
  CANR1X1 U1387 ( .A(n288), .B(n1610), .C(n283), .Z(n281) );
  CENX1 U1388 ( .A(n1649), .B(n1634), .Z(n1423) );
  CANR1XL U1389 ( .A(n373), .B(n1617), .C(n370), .Z(n368) );
  CIVX3 U1390 ( .A(n1692), .Z(n1691) );
  CANR1X1 U1391 ( .A(n312), .B(n293), .C(n294), .Z(n292) );
  CNR2X1 U1392 ( .A(n295), .B(n298), .Z(n293) );
  CIVX2 U1393 ( .A(n30), .Z(n1679) );
  CIVX2 U1394 ( .A(n39), .Z(n1685) );
  CAOR1XL U1395 ( .A(n312), .B(n293), .C(n294), .Z(n1560) );
  CNIVX2 U1396 ( .A(n124), .Z(n1561) );
  CNIVX2 U1397 ( .A(n122), .Z(n1562) );
  CNIVX2 U1398 ( .A(n126), .Z(n1563) );
  CIVX2 U1399 ( .A(n21), .Z(n1673) );
  CNIVX2 U1400 ( .A(n128), .Z(n1564) );
  CIVX2 U1401 ( .A(n1646), .Z(n1585) );
  COR2X1 U1402 ( .A(n1136), .B(n865), .Z(n1565) );
  CIVX1 U1403 ( .A(n1688), .Z(n1566) );
  CEOXL U1404 ( .A(n236), .B(n1567), .Z(product[26]) );
  CND2X1 U1405 ( .A(n389), .B(n235), .Z(n1567) );
  CFA1XL U1406 ( .A(n940), .B(n870), .CI(n1000), .CO(n478), .S(n479) );
  COND2XL U1407 ( .A(n61), .B(n1238), .C(n1237), .D(n1631), .Z(n957) );
  CENX1 U1408 ( .A(n1653), .B(b[25]), .Z(n1398) );
  CFA1XL U1409 ( .A(n961), .B(n1081), .CI(n1053), .CO(n554), .S(n555) );
  CND2X1 U1410 ( .A(n216), .B(n228), .Z(n214) );
  CENXL U1411 ( .A(n220), .B(n1568), .Z(product[28]) );
  CAN2XL U1412 ( .A(n387), .B(n219), .Z(n1568) );
  CENXL U1413 ( .A(n227), .B(n1569), .Z(product[27]) );
  CAN2X1 U1414 ( .A(n388), .B(n226), .Z(n1569) );
  CENXL U1415 ( .A(n1651), .B(n1647), .Z(n1169) );
  CENXL U1416 ( .A(n1563), .B(n1647), .Z(n1166) );
  CIVXL U1417 ( .A(n1644), .Z(n1475) );
  CENX2 U1418 ( .A(n1682), .B(a[10]), .Z(n50) );
  COND2XL U1419 ( .A(n44), .B(n1686), .C(n42), .D(n1304), .Z(n861) );
  CIVX1 U1420 ( .A(n279), .Z(n278) );
  CIVX3 U1421 ( .A(n1689), .Z(n1687) );
  CENX1 U1422 ( .A(n1687), .B(n1652), .Z(n1277) );
  CENXL U1423 ( .A(n1649), .B(n1684), .Z(n1303) );
  CENX1 U1424 ( .A(n1649), .B(n109), .Z(n1143) );
  CENXL U1425 ( .A(n1649), .B(n1647), .Z(n1170) );
  CENX1 U1426 ( .A(n1649), .B(n104), .Z(n1150) );
  CIVX4 U1427 ( .A(n1570), .Z(n1688) );
  CENX2 U1428 ( .A(n1682), .B(a[10]), .Z(n1597) );
  CIVX2 U1429 ( .A(n48), .Z(n1570) );
  CIVX2 U1430 ( .A(n48), .Z(n1689) );
  CNR2IX1 U1431 ( .B(n1559), .A(n1631), .Z(n975) );
  CIVX1 U1432 ( .A(n330), .Z(n329) );
  CND2IXL U1433 ( .B(n1559), .A(n1691), .Z(n1256) );
  CNR2X1 U1434 ( .A(n487), .B(n512), .Z(n1571) );
  CNR2XL U1435 ( .A(n487), .B(n512), .Z(n1572) );
  CNR2XL U1436 ( .A(n487), .B(n512), .Z(n218) );
  CENX4 U1437 ( .A(n1644), .B(a[18]), .Z(n82) );
  COND2X1 U1438 ( .A(n85), .B(n1187), .C(n1186), .D(n82), .Z(n909) );
  CND2IX2 U1439 ( .B(n1603), .A(n50), .Z(n53) );
  CEOX2 U1440 ( .A(n1693), .B(a[16]), .Z(n1573) );
  CEOX1 U1441 ( .A(n1693), .B(a[16]), .Z(n1625) );
  CNIVX1 U1442 ( .A(n1062), .Z(n1574) );
  CENXL U1443 ( .A(n1644), .B(n146), .Z(n1201) );
  COND2XL U1444 ( .A(n36), .B(n1306), .C(n1305), .D(n33), .Z(n1022) );
  COND2XL U1445 ( .A(n36), .B(n1308), .C(n1307), .D(n33), .Z(n1024) );
  COND2XL U1446 ( .A(n36), .B(n1307), .C(n1306), .D(n33), .Z(n1023) );
  COND2XL U1447 ( .A(n36), .B(n1322), .C(n1321), .D(n33), .Z(n1038) );
  COND2XL U1448 ( .A(n36), .B(n1678), .C(n33), .D(n1331), .Z(n862) );
  COND2XL U1449 ( .A(n36), .B(n1326), .C(n1325), .D(n33), .Z(n1042) );
  COND2XL U1450 ( .A(n1330), .B(n36), .C(n1329), .D(n33), .Z(n1046) );
  COND2XL U1451 ( .A(n36), .B(n1323), .C(n1322), .D(n33), .Z(n1039) );
  COND2XL U1452 ( .A(n36), .B(n1309), .C(n1308), .D(n33), .Z(n1025) );
  COND2XL U1453 ( .A(n36), .B(n1318), .C(n1317), .D(n33), .Z(n1034) );
  COND2XL U1454 ( .A(n36), .B(n1316), .C(n1315), .D(n33), .Z(n1032) );
  COND2XL U1455 ( .A(n36), .B(n1314), .C(n1313), .D(n33), .Z(n1030) );
  CIVX2 U1456 ( .A(n1623), .Z(n1629) );
  CANR1X1 U1457 ( .A(n229), .B(n216), .C(n217), .Z(n1575) );
  CANR1XL U1458 ( .A(n229), .B(n216), .C(n217), .Z(n215) );
  CENXL U1459 ( .A(n208), .B(n1576), .Z(product[30]) );
  CAN2XL U1460 ( .A(n385), .B(n207), .Z(n1576) );
  COND1X2 U1461 ( .A(n240), .B(n234), .C(n235), .Z(n229) );
  CND2X1 U1462 ( .A(n563), .B(n586), .Z(n240) );
  CENX1 U1463 ( .A(n1674), .B(n153), .Z(n1311) );
  COND1X1 U1464 ( .A(n330), .B(n313), .C(n314), .Z(n312) );
  CND2XL U1465 ( .A(n320), .B(n1612), .Z(n313) );
  COND2X1 U1466 ( .A(n77), .B(n1209), .C(n1208), .D(n1635), .Z(n930) );
  CFA1XL U1467 ( .A(n851), .B(n924), .CI(n978), .CO(n480), .S(n481) );
  COND2X1 U1468 ( .A(n77), .B(n1202), .C(n1201), .D(n1635), .Z(n923) );
  COND1XL U1469 ( .A(n214), .B(n242), .C(n215), .Z(n213) );
  CENX2 U1470 ( .A(n1646), .B(a[22]), .Z(n95) );
  CEOX1 U1471 ( .A(a[22]), .B(n1647), .Z(n1447) );
  CENXL U1472 ( .A(n1659), .B(n130), .Z(n1384) );
  CENXL U1473 ( .A(n1690), .B(n130), .Z(n1249) );
  CENXL U1474 ( .A(n130), .B(n1647), .Z(n1164) );
  CANR1X1 U1475 ( .A(n1612), .B(n321), .C(n316), .Z(n314) );
  CNR2X1 U1476 ( .A(n234), .B(n239), .Z(n228) );
  CENXL U1477 ( .A(n1653), .B(b[30]), .Z(n1393) );
  CENXL U1478 ( .A(n1653), .B(b[29]), .Z(n1394) );
  CENXL U1479 ( .A(n1653), .B(n132), .Z(n1416) );
  CENXL U1480 ( .A(n1653), .B(b[28]), .Z(n1395) );
  CENXL U1481 ( .A(n1653), .B(b[27]), .Z(n1396) );
  CENXL U1482 ( .A(n1653), .B(n155), .Z(n1402) );
  CENXL U1483 ( .A(n1653), .B(n156), .Z(n1401) );
  CENXL U1484 ( .A(n1653), .B(n154), .Z(n1403) );
  COND2X1 U1485 ( .A(n77), .B(n1210), .C(n1209), .D(n1635), .Z(n931) );
  CENXL U1486 ( .A(n1687), .B(n155), .Z(n1257) );
  CENXL U1487 ( .A(n1687), .B(n1564), .Z(n1273) );
  CENXL U1488 ( .A(n1687), .B(n153), .Z(n1259) );
  CENXL U1489 ( .A(n1687), .B(n1563), .Z(n1274) );
  CENXL U1490 ( .A(n1687), .B(n154), .Z(n1258) );
  CENXL U1491 ( .A(n1687), .B(n1561), .Z(n1275) );
  CENXL U1492 ( .A(n1687), .B(n1562), .Z(n1276) );
  COND2XL U1493 ( .A(n77), .B(n1201), .C(n1200), .D(n1635), .Z(n922) );
  COND2XL U1494 ( .A(n77), .B(n1204), .C(n1203), .D(n1635), .Z(n925) );
  COND2XL U1495 ( .A(n1215), .B(n77), .C(n1635), .D(n1214), .Z(n936) );
  COND2XL U1496 ( .A(n77), .B(n1203), .C(n1202), .D(n1635), .Z(n924) );
  COND2XL U1497 ( .A(n77), .B(n1213), .C(n1212), .D(n1635), .Z(n934) );
  CENXL U1498 ( .A(n1688), .B(n138), .Z(n1268) );
  CND2IXL U1499 ( .B(n1559), .A(n1688), .Z(n1279) );
  CENXL U1500 ( .A(n1649), .B(n1688), .Z(n1278) );
  CENXL U1501 ( .A(n1688), .B(n136), .Z(n1269) );
  CENXL U1502 ( .A(n1688), .B(n152), .Z(n1260) );
  CENXL U1503 ( .A(n1688), .B(n142), .Z(n1266) );
  CENXL U1504 ( .A(n1688), .B(n146), .Z(n1264) );
  CENXL U1505 ( .A(n1688), .B(n148), .Z(n1263) );
  CENXL U1506 ( .A(n1688), .B(n151), .Z(n1261) );
  CENX2 U1507 ( .A(a[10]), .B(n1688), .Z(n1603) );
  CANR1X1 U1508 ( .A(n1607), .B(n1577), .C(n210), .Z(n208) );
  CANR1X1 U1509 ( .A(n1606), .B(n1557), .C(n1605), .Z(n199) );
  CND2X2 U1510 ( .A(n95), .B(n1447), .Z(n97) );
  CEO3X1 U1511 ( .A(n662), .B(n647), .C(n649), .Z(n639) );
  CND2X1 U1512 ( .A(n662), .B(n647), .Z(n1578) );
  CND2X1 U1513 ( .A(n662), .B(n649), .Z(n1579) );
  CND2X1 U1514 ( .A(n647), .B(n649), .Z(n1580) );
  CEOX1 U1515 ( .A(n636), .B(n619), .Z(n1581) );
  CND2X1 U1516 ( .A(n636), .B(n619), .Z(n1582) );
  CND2X1 U1517 ( .A(n636), .B(n638), .Z(n1583) );
  CND2X1 U1518 ( .A(n619), .B(n638), .Z(n1584) );
  CND2X1 U1519 ( .A(a[20]), .B(n1585), .Z(n1586) );
  CND2XL U1520 ( .A(n1594), .B(n1646), .Z(n1587) );
  CND2X1 U1521 ( .A(n1586), .B(n1587), .Z(n1448) );
  CHA1XL U1522 ( .A(n930), .B(n904), .CO(n628), .S(n629) );
  CENXL U1523 ( .A(n1695), .B(n140), .Z(n1223) );
  CENXL U1524 ( .A(n1644), .B(n140), .Z(n1204) );
  CENXL U1525 ( .A(n1645), .B(n144), .Z(n1185) );
  CENXL U1526 ( .A(n1676), .B(n144), .Z(n1317) );
  CENXL U1527 ( .A(n1663), .B(n144), .Z(n1377) );
  CENXL U1528 ( .A(n1644), .B(n144), .Z(n1202) );
  CENXL U1529 ( .A(n1634), .B(n144), .Z(n1410) );
  CENXL U1530 ( .A(n1683), .B(n144), .Z(n1290) );
  CENXL U1531 ( .A(n1670), .B(n144), .Z(n1346) );
  CENXL U1532 ( .A(n1687), .B(n144), .Z(n1265) );
  COND2X1 U1533 ( .A(n91), .B(n1177), .C(n1176), .D(n89), .Z(n900) );
  CNIVX4 U1534 ( .A(n79), .Z(n1645) );
  COND2X1 U1535 ( .A(n1198), .B(n85), .C(n82), .D(n1197), .Z(n920) );
  CENXL U1536 ( .A(n1676), .B(b[25]), .Z(n1305) );
  CENXL U1537 ( .A(n1666), .B(b[25]), .Z(n1334) );
  CENXL U1538 ( .A(n1658), .B(b[25]), .Z(n1365) );
  CND2X2 U1539 ( .A(n1449), .B(n82), .Z(n85) );
  COND1X1 U1540 ( .A(n352), .B(n340), .C(n341), .Z(n339) );
  CANR1X1 U1541 ( .A(n1615), .B(n357), .C(n354), .Z(n352) );
  CIVXL U1542 ( .A(n889), .Z(n1588) );
  CIVX2 U1543 ( .A(n1588), .Z(n1589) );
  COND2XL U1544 ( .A(n97), .B(n1164), .C(n1163), .D(n95), .Z(n888) );
  COND2XL U1545 ( .A(n97), .B(n1165), .C(n1164), .D(n95), .Z(n889) );
  COND2XL U1546 ( .A(n1170), .B(n97), .C(n95), .D(n1169), .Z(n894) );
  COND2XL U1547 ( .A(n97), .B(n1166), .C(n95), .D(n1165), .Z(n890) );
  CNR2IXL U1548 ( .B(n1559), .A(n95), .Z(n895) );
  COND2X1 U1549 ( .A(n1171), .B(n95), .C(n1472), .D(n97), .Z(n854) );
  CENXL U1550 ( .A(n1690), .B(n134), .Z(n1247) );
  CENXL U1551 ( .A(n1687), .B(n134), .Z(n1270) );
  CENXL U1552 ( .A(n134), .B(n1647), .Z(n1162) );
  CENXL U1553 ( .A(n1645), .B(n134), .Z(n1190) );
  CEOX2 U1554 ( .A(a[6]), .B(n1677), .Z(n1455) );
  CIVXL U1555 ( .A(n39), .Z(n1686) );
  CIVX2 U1556 ( .A(n100), .Z(n1590) );
  CIVX2 U1557 ( .A(n1590), .Z(n1591) );
  CIVX2 U1558 ( .A(n1590), .Z(n1592) );
  CND2IXL U1559 ( .B(n1559), .A(n109), .Z(n1144) );
  CND2X2 U1560 ( .A(n1645), .B(a[20]), .Z(n1595) );
  CND2X2 U1561 ( .A(n1593), .B(n1594), .Z(n1596) );
  CND2X4 U1562 ( .A(n1595), .B(n1596), .Z(n89) );
  CIVX1 U1563 ( .A(n1645), .Z(n1593) );
  CIVX2 U1564 ( .A(a[20]), .Z(n1594) );
  COND2X1 U1565 ( .A(n91), .B(n1175), .C(n1174), .D(n89), .Z(n898) );
  COND2X1 U1566 ( .A(n91), .B(n1176), .C(n1175), .D(n89), .Z(n899) );
  COND2X1 U1567 ( .A(n91), .B(n1174), .C(n1173), .D(n89), .Z(n897) );
  COND2X1 U1568 ( .A(n1183), .B(n91), .C(n89), .D(n1182), .Z(n906) );
  COND2XL U1569 ( .A(n91), .B(n1181), .C(n89), .D(n1180), .Z(n904) );
  CIVX3 U1570 ( .A(n1685), .Z(n1682) );
  COND1X1 U1571 ( .A(n299), .B(n295), .C(n296), .Z(n294) );
  COR2XL U1572 ( .A(n53), .B(n1272), .Z(n1598) );
  COR2XL U1573 ( .A(n1271), .B(n1597), .Z(n1599) );
  CND2X1 U1574 ( .A(n1598), .B(n1599), .Z(n990) );
  CENXL U1575 ( .A(n1687), .B(n132), .Z(n1271) );
  COR2XL U1576 ( .A(n53), .B(n1277), .Z(n1600) );
  COR2XL U1577 ( .A(n1276), .B(n1597), .Z(n1601) );
  CND2X1 U1578 ( .A(n1600), .B(n1601), .Z(n995) );
  COND2X1 U1579 ( .A(n44), .B(n1287), .C(n1286), .D(n42), .Z(n1004) );
  CND2X1 U1580 ( .A(n1610), .B(n1611), .Z(n280) );
  CNIVX1 U1581 ( .A(n1655), .Z(n1634) );
  CIVX1 U1582 ( .A(n1656), .Z(n1653) );
  COND2X1 U1583 ( .A(n9), .B(n1399), .C(n6), .D(n1398), .Z(n1112) );
  CNR2IX1 U1584 ( .B(n1559), .A(n33), .Z(n1047) );
  CANR1XL U1585 ( .A(n365), .B(n1618), .C(n362), .Z(n360) );
  CANR1XL U1586 ( .A(n381), .B(n1619), .C(n378), .Z(n376) );
  CND2XL U1587 ( .A(n412), .B(n375), .Z(n194) );
  CEO3X1 U1588 ( .A(n452), .B(n450), .C(n448), .Z(n422) );
  COND2XL U1589 ( .A(n18), .B(n1389), .C(n15), .D(n1388), .Z(n1103) );
  CNR2IXL U1590 ( .B(n1559), .A(n24), .Z(n1075) );
  CENX1 U1591 ( .A(n1684), .B(n153), .Z(n1284) );
  CENX1 U1592 ( .A(n1671), .B(n152), .Z(n1341) );
  CENX1 U1593 ( .A(n1658), .B(n156), .Z(n1368) );
  CEOX2 U1594 ( .A(n1661), .B(a[4]), .Z(n1624) );
  CIVX4 U1595 ( .A(n1624), .Z(n24) );
  CENX2 U1596 ( .A(n1648), .B(a[26]), .Z(n105) );
  CIVX2 U1597 ( .A(n1655), .Z(n1621) );
  CENX2 U1598 ( .A(a[0]), .B(n1621), .Z(n1458) );
  CENX1 U1599 ( .A(n1676), .B(n150), .Z(n1314) );
  CENX1 U1600 ( .A(n1671), .B(n150), .Z(n1343) );
  CENX1 U1601 ( .A(n1634), .B(n150), .Z(n1407) );
  CENX1 U1602 ( .A(n1664), .B(n150), .Z(n1374) );
  CENX1 U1603 ( .A(n1684), .B(n150), .Z(n1287) );
  CENXL U1604 ( .A(n1688), .B(n150), .Z(n1262) );
  CANR1X1 U1605 ( .A(n308), .B(n1608), .C(n301), .Z(n299) );
  CIVX1 U1606 ( .A(n306), .Z(n308) );
  CEOXL U1607 ( .A(n177), .B(n286), .Z(product[20]) );
  CND2XL U1608 ( .A(n1610), .B(n285), .Z(n177) );
  CEOXL U1609 ( .A(n176), .B(n278), .Z(product[21]) );
  CND2XL U1610 ( .A(n394), .B(n273), .Z(n176) );
  CND2XL U1611 ( .A(n1612), .B(n318), .Z(n182) );
  CEOXL U1612 ( .A(n181), .B(n311), .Z(product[16]) );
  CND2XL U1613 ( .A(n399), .B(n306), .Z(n181) );
  CND2XL U1614 ( .A(n1611), .B(n290), .Z(n178) );
  CND2XL U1615 ( .A(n1608), .B(n303), .Z(n180) );
  CND2XL U1616 ( .A(n399), .B(n1608), .Z(n298) );
  CND2XL U1617 ( .A(n587), .B(n608), .Z(n250) );
  CANR1X1 U1618 ( .A(n275), .B(n1609), .C(n268), .Z(n262) );
  CIVX1 U1619 ( .A(n273), .Z(n275) );
  CIVXL U1620 ( .A(n262), .Z(n264) );
  CANR1X1 U1621 ( .A(n331), .B(n339), .C(n332), .Z(n330) );
  CNR2XL U1622 ( .A(n333), .B(n336), .Z(n331) );
  CENX1 U1623 ( .A(n1602), .B(n633), .Z(n631) );
  CENX1 U1624 ( .A(n635), .B(n652), .Z(n1602) );
  CNR2XL U1625 ( .A(n322), .B(n327), .Z(n320) );
  CND2XL U1626 ( .A(n1614), .B(n345), .Z(n187) );
  CND2XL U1627 ( .A(n404), .B(n337), .Z(n186) );
  CND2XL U1628 ( .A(n1615), .B(n356), .Z(n189) );
  CND2XL U1629 ( .A(n1613), .B(n350), .Z(n188) );
  CND2XL U1630 ( .A(n402), .B(n328), .Z(n184) );
  CND2XL U1631 ( .A(n707), .B(n722), .Z(n296) );
  CND2XL U1632 ( .A(n767), .B(n778), .Z(n323) );
  COND1X1 U1633 ( .A(n358), .B(n360), .C(n359), .Z(n357) );
  CND2XL U1634 ( .A(n430), .B(n415), .Z(n198) );
  CND2XL U1635 ( .A(n791), .B(n800), .Z(n334) );
  CND2XL U1636 ( .A(n408), .B(n359), .Z(n190) );
  CND2IXL U1637 ( .B(n366), .A(n367), .Z(n192) );
  CND2XL U1638 ( .A(n1617), .B(n372), .Z(n193) );
  CND2XL U1639 ( .A(n1618), .B(n364), .Z(n191) );
  CEOXL U1640 ( .A(n376), .B(n194), .Z(product[3]) );
  CND2XL U1641 ( .A(n1619), .B(n380), .Z(n195) );
  CND2XL U1642 ( .A(n843), .B(n846), .Z(n367) );
  CND2XL U1643 ( .A(n849), .B(n1104), .Z(n375) );
  CEO3X1 U1644 ( .A(n434), .B(n416), .C(n432), .Z(n415) );
  CEO3X1 U1645 ( .A(n436), .B(n418), .C(n417), .Z(n416) );
  CEO3X1 U1646 ( .A(n420), .B(n438), .C(n419), .Z(n417) );
  CAN2XL U1647 ( .A(n1565), .B(n383), .Z(product[1]) );
  CIVX2 U1648 ( .A(n1680), .Z(n1677) );
  COND2XL U1649 ( .A(n36), .B(n1313), .C(n1312), .D(n33), .Z(n1029) );
  CNR2IXL U1650 ( .B(n1559), .A(n42), .Z(n1021) );
  COND2XL U1651 ( .A(n36), .B(n1329), .C(n1328), .D(n33), .Z(n1045) );
  COND2XL U1652 ( .A(n97), .B(n1162), .C(n1161), .D(n95), .Z(n886) );
  CNR2IXL U1653 ( .B(n1559), .A(n6), .Z(product[0]) );
  COR2X2 U1654 ( .A(n1622), .B(n1573), .Z(n77) );
  CENX1 U1655 ( .A(n1644), .B(a[16]), .Z(n1622) );
  CENX1 U1656 ( .A(n1667), .B(n155), .Z(n1338) );
  CND2X2 U1657 ( .A(n1591), .B(n1446), .Z(n102) );
  CEOX1 U1658 ( .A(a[24]), .B(n1648), .Z(n1446) );
  CENXL U1659 ( .A(n1684), .B(n157), .Z(n1280) );
  CNIVX1 U1660 ( .A(n116), .Z(n1649) );
  CENXL U1661 ( .A(n1695), .B(n142), .Z(n1222) );
  CENXL U1662 ( .A(n1690), .B(n140), .Z(n1244) );
  CENXL U1663 ( .A(n1691), .B(n144), .Z(n1242) );
  CENXL U1664 ( .A(n1696), .B(n144), .Z(n1221) );
  CNIVX4 U1665 ( .A(n71), .Z(n1644) );
  CNIVX2 U1666 ( .A(n120), .Z(n1651) );
  CND2XL U1667 ( .A(n1443), .B(n114), .Z(n115) );
  CANR1XL U1668 ( .A(n390), .B(n241), .C(n238), .Z(n236) );
  CEOXL U1669 ( .A(n213), .B(n1604), .Z(product[29]) );
  CAN2XL U1670 ( .A(n1607), .B(n212), .Z(n1604) );
  CENX1 U1671 ( .A(n251), .B(n173), .Z(product[24]) );
  COND1XL U1672 ( .A(n252), .B(n278), .C(n253), .Z(n251) );
  CND2XL U1673 ( .A(n263), .B(n392), .Z(n252) );
  CENX1 U1674 ( .A(n241), .B(n172), .Z(product[25]) );
  COND1XL U1675 ( .A(n223), .B(n231), .C(n226), .Z(n222) );
  CANR1XL U1676 ( .A(n228), .B(n241), .C(n229), .Z(n227) );
  CANR1XL U1677 ( .A(n221), .B(n241), .C(n222), .Z(n220) );
  CNR2IXL U1678 ( .B(n228), .A(n223), .Z(n221) );
  CAOR1X1 U1679 ( .A(n210), .B(n385), .C(n205), .Z(n1605) );
  CAN2XL U1680 ( .A(n385), .B(n1607), .Z(n1606) );
  CANR1XL U1681 ( .A(n392), .B(n264), .C(n257), .Z(n253) );
  CENX1 U1682 ( .A(n304), .B(n180), .Z(product[17]) );
  COND1XL U1683 ( .A(n305), .B(n311), .C(n306), .Z(n304) );
  CENX1 U1684 ( .A(n297), .B(n179), .Z(product[18]) );
  CND2X1 U1685 ( .A(n397), .B(n296), .Z(n179) );
  COND1XL U1686 ( .A(n298), .B(n311), .C(n299), .Z(n297) );
  CENX1 U1687 ( .A(n271), .B(n175), .Z(product[22]) );
  CND2X1 U1688 ( .A(n1609), .B(n270), .Z(n175) );
  COND1XL U1689 ( .A(n272), .B(n278), .C(n273), .Z(n271) );
  CENX1 U1690 ( .A(n260), .B(n174), .Z(product[23]) );
  CND2XL U1691 ( .A(n392), .B(n259), .Z(n174) );
  COND1XL U1692 ( .A(n261), .B(n278), .C(n262), .Z(n260) );
  CENX1 U1693 ( .A(n1560), .B(n178), .Z(product[19]) );
  CNR2X1 U1694 ( .A(n563), .B(n586), .Z(n239) );
  CANR1XL U1695 ( .A(n1611), .B(n1560), .C(n288), .Z(n286) );
  CEOX1 U1696 ( .A(n183), .B(n324), .Z(product[14]) );
  CND2X1 U1697 ( .A(n401), .B(n323), .Z(n183) );
  CANR1XL U1698 ( .A(n402), .B(n329), .C(n326), .Z(n324) );
  CEOX1 U1699 ( .A(n182), .B(n319), .Z(product[15]) );
  CANR1XL U1700 ( .A(n320), .B(n329), .C(n321), .Z(n319) );
  COR2X1 U1701 ( .A(n459), .B(n486), .Z(n1607) );
  CNR2X1 U1702 ( .A(n587), .B(n608), .Z(n249) );
  CND2X1 U1703 ( .A(n513), .B(n538), .Z(n226) );
  CND2X1 U1704 ( .A(n1609), .B(n394), .Z(n261) );
  CND2X1 U1705 ( .A(n539), .B(n562), .Z(n235) );
  CND2X1 U1706 ( .A(n487), .B(n512), .Z(n219) );
  CND2X1 U1707 ( .A(n1614), .B(n1613), .Z(n340) );
  CNR2X1 U1708 ( .A(n707), .B(n722), .Z(n295) );
  COND1XL U1709 ( .A(n337), .B(n333), .C(n334), .Z(n332) );
  COND1XL U1710 ( .A(n328), .B(n322), .C(n323), .Z(n321) );
  CNR2X1 U1711 ( .A(n767), .B(n778), .Z(n322) );
  CENX1 U1712 ( .A(n188), .B(n351), .Z(product[9]) );
  CENX1 U1713 ( .A(n335), .B(n185), .Z(product[12]) );
  CND2X1 U1714 ( .A(n403), .B(n334), .Z(n185) );
  COND1XL U1715 ( .A(n336), .B(n338), .C(n337), .Z(n335) );
  CENX1 U1716 ( .A(n329), .B(n184), .Z(product[13]) );
  CNR2X1 U1717 ( .A(n739), .B(n752), .Z(n305) );
  COR2X1 U1718 ( .A(n723), .B(n738), .Z(n1608) );
  CEOX1 U1719 ( .A(n346), .B(n187), .Z(product[10]) );
  CANR1XL U1720 ( .A(n1613), .B(n351), .C(n348), .Z(n346) );
  CEOX1 U1721 ( .A(n186), .B(n338), .Z(product[11]) );
  COR2X1 U1722 ( .A(n631), .B(n650), .Z(n1609) );
  COR2X1 U1723 ( .A(n671), .B(n688), .Z(n1610) );
  COR2X1 U1724 ( .A(n689), .B(n706), .Z(n1611) );
  COR2X1 U1725 ( .A(n753), .B(n766), .Z(n1612) );
  CND2X1 U1726 ( .A(n651), .B(n670), .Z(n273) );
  CND2X1 U1727 ( .A(n739), .B(n752), .Z(n306) );
  CND2X1 U1728 ( .A(n1638), .B(n630), .Z(n259) );
  CND2X1 U1729 ( .A(n689), .B(n706), .Z(n290) );
  CND2X1 U1730 ( .A(n631), .B(n650), .Z(n270) );
  CND2X1 U1731 ( .A(n671), .B(n688), .Z(n285) );
  CND2X1 U1732 ( .A(n753), .B(n766), .Z(n318) );
  CND2X1 U1733 ( .A(n723), .B(n738), .Z(n303) );
  COND1XL U1734 ( .A(n376), .B(n374), .C(n375), .Z(n373) );
  CND2X1 U1735 ( .A(n1616), .B(n198), .Z(n166) );
  CNR2X1 U1736 ( .A(n801), .B(n810), .Z(n336) );
  CNR2X1 U1737 ( .A(n791), .B(n800), .Z(n333) );
  CNR2X1 U1738 ( .A(n779), .B(n790), .Z(n327) );
  COR2X1 U1739 ( .A(n819), .B(n826), .Z(n1613) );
  COR2X1 U1740 ( .A(n811), .B(n818), .Z(n1614) );
  CND2X1 U1741 ( .A(n779), .B(n790), .Z(n328) );
  CND2X1 U1742 ( .A(n801), .B(n810), .Z(n337) );
  CND2X1 U1743 ( .A(n819), .B(n826), .Z(n350) );
  CND2X1 U1744 ( .A(n827), .B(n832), .Z(n356) );
  CND2X1 U1745 ( .A(n811), .B(n818), .Z(n345) );
  COR2X1 U1746 ( .A(n827), .B(n832), .Z(n1615) );
  COR2X1 U1747 ( .A(n430), .B(n415), .Z(n1616) );
  CENX1 U1748 ( .A(n193), .B(n373), .Z(product[4]) );
  CENX1 U1749 ( .A(n191), .B(n365), .Z(product[6]) );
  CEOXL U1750 ( .A(n360), .B(n190), .Z(product[7]) );
  CENX1 U1751 ( .A(n195), .B(n381), .Z(product[2]) );
  CNR2X1 U1752 ( .A(n843), .B(n846), .Z(n366) );
  CNR2X1 U1753 ( .A(n833), .B(n838), .Z(n358) );
  CNR2X1 U1754 ( .A(n849), .B(n1104), .Z(n374) );
  COR2X1 U1755 ( .A(n847), .B(n848), .Z(n1617) );
  COR2X1 U1756 ( .A(n839), .B(n842), .Z(n1618) );
  CND2X1 U1757 ( .A(n1135), .B(n1105), .Z(n380) );
  CND2X1 U1758 ( .A(n847), .B(n848), .Z(n372) );
  CND2X1 U1759 ( .A(n839), .B(n842), .Z(n364) );
  CND2X1 U1760 ( .A(n833), .B(n838), .Z(n359) );
  COR2X1 U1761 ( .A(n1135), .B(n1105), .Z(n1619) );
  CENX1 U1762 ( .A(n1675), .B(n1562), .Z(n1328) );
  CENX1 U1763 ( .A(n1675), .B(n1564), .Z(n1325) );
  CENX1 U1764 ( .A(n1681), .B(n1563), .Z(n1299) );
  CENX1 U1765 ( .A(n1681), .B(n1564), .Z(n1298) );
  CENX1 U1766 ( .A(n1675), .B(n1563), .Z(n1326) );
  CENX1 U1767 ( .A(n1675), .B(n1561), .Z(n1327) );
  CENX1 U1768 ( .A(n1693), .B(n1564), .Z(n1229) );
  CENX1 U1769 ( .A(n1562), .B(n1645), .Z(n1196) );
  CENX1 U1770 ( .A(n1654), .B(n1564), .Z(n1418) );
  CENX1 U1771 ( .A(n1654), .B(n1651), .Z(n1422) );
  CENX1 U1772 ( .A(n1654), .B(n1562), .Z(n1421) );
  CENX1 U1773 ( .A(n1654), .B(n1563), .Z(n1419) );
  CENX1 U1774 ( .A(n1654), .B(n1561), .Z(n1420) );
  CNR2IX1 U1775 ( .B(n1559), .A(n110), .Z(n871) );
  CENX1 U1776 ( .A(n1651), .B(n1645), .Z(n1197) );
  CENX1 U1777 ( .A(n1668), .B(n1563), .Z(n1355) );
  CENX1 U1778 ( .A(n1669), .B(n1562), .Z(n1357) );
  CENX1 U1779 ( .A(n1669), .B(n1561), .Z(n1356) );
  CNR2IXL U1780 ( .B(n1559), .A(n15), .Z(n1105) );
  CENX1 U1781 ( .A(n1564), .B(n1646), .Z(n1178) );
  CENX1 U1782 ( .A(n1690), .B(n1651), .Z(n1254) );
  CENX1 U1783 ( .A(n1682), .B(n1652), .Z(n1302) );
  CENX1 U1784 ( .A(n1682), .B(n1562), .Z(n1301) );
  CENX1 U1785 ( .A(n1690), .B(n1563), .Z(n1251) );
  CENX1 U1786 ( .A(n1690), .B(n1564), .Z(n1250) );
  CENX1 U1787 ( .A(n1690), .B(n1561), .Z(n1252) );
  CENX1 U1788 ( .A(n1690), .B(n1562), .Z(n1253) );
  CENX1 U1789 ( .A(n1675), .B(n1651), .Z(n1329) );
  CENX1 U1790 ( .A(n1651), .B(n1648), .Z(n1158) );
  CENX1 U1791 ( .A(n1562), .B(n1648), .Z(n1157) );
  CENX1 U1792 ( .A(n1564), .B(n1647), .Z(n1165) );
  CENX1 U1793 ( .A(n1561), .B(n1648), .Z(n1156) );
  CENX1 U1794 ( .A(n1561), .B(n1647), .Z(n1167) );
  CENX1 U1795 ( .A(n1564), .B(n1648), .Z(n1154) );
  CENX1 U1796 ( .A(n1562), .B(n1646), .Z(n1181) );
  CENX1 U1797 ( .A(n1562), .B(n1647), .Z(n1168) );
  CENX1 U1798 ( .A(n1563), .B(n1648), .Z(n1155) );
  CENX1 U1799 ( .A(n1694), .B(n1562), .Z(n1232) );
  CENX1 U1800 ( .A(n1563), .B(n1646), .Z(n1179) );
  CENX1 U1801 ( .A(n1651), .B(n1646), .Z(n1182) );
  CENX1 U1802 ( .A(n1561), .B(n1646), .Z(n1180) );
  CENX1 U1803 ( .A(n1649), .B(n1677), .Z(n1330) );
  CENX1 U1804 ( .A(n1649), .B(n1648), .Z(n1159) );
  CENX1 U1805 ( .A(n1694), .B(n1561), .Z(n1231) );
  CENX1 U1806 ( .A(n1660), .B(n1561), .Z(n1387) );
  CENX1 U1807 ( .A(n1661), .B(n1651), .Z(n1389) );
  CENX1 U1808 ( .A(n1660), .B(n1564), .Z(n1385) );
  CENX1 U1809 ( .A(n1660), .B(n1563), .Z(n1386) );
  CENX1 U1810 ( .A(n1649), .B(n1646), .Z(n1183) );
  CENX1 U1811 ( .A(n1649), .B(n1672), .Z(n1359) );
  CNR2IX1 U1812 ( .B(n1559), .A(n114), .Z(n867) );
  CNR2IX1 U1813 ( .B(n1559), .A(n1635), .Z(n937) );
  CNR2IX1 U1814 ( .B(n1559), .A(n105), .Z(n877) );
  CIVX8 U1815 ( .A(n1692), .Z(n1690) );
  CNIVX1 U1816 ( .A(n915), .Z(n1633) );
  CNR2IX1 U1817 ( .B(n1559), .A(n1592), .Z(n885) );
  CEOX1 U1818 ( .A(n872), .B(n886), .Z(n429) );
  CIVXL U1819 ( .A(n1698), .Z(n1695) );
  CENX1 U1820 ( .A(n1669), .B(b[27]), .Z(n1332) );
  CENX1 U1821 ( .A(n1695), .B(n138), .Z(n1224) );
  CENX1 U1822 ( .A(n1667), .B(n154), .Z(n1339) );
  CENX1 U1823 ( .A(n1695), .B(n132), .Z(n1227) );
  CENX1 U1824 ( .A(n1676), .B(n156), .Z(n1308) );
  CENX1 U1825 ( .A(n1690), .B(n138), .Z(n1245) );
  CENX1 U1826 ( .A(n1671), .B(n148), .Z(n1344) );
  CENX1 U1827 ( .A(n1676), .B(n142), .Z(n1318) );
  CENX1 U1828 ( .A(n1684), .B(n136), .Z(n1294) );
  CENX1 U1829 ( .A(n1671), .B(n151), .Z(n1342) );
  CENX1 U1830 ( .A(n1690), .B(n136), .Z(n1246) );
  CENX1 U1831 ( .A(n1684), .B(n148), .Z(n1288) );
  CENX1 U1832 ( .A(n1684), .B(n154), .Z(n1283) );
  CENX1 U1833 ( .A(n1684), .B(n155), .Z(n1282) );
  CENX1 U1834 ( .A(n1676), .B(n136), .Z(n1321) );
  CENX1 U1835 ( .A(n1694), .B(n136), .Z(n1225) );
  CENX1 U1836 ( .A(n1683), .B(n138), .Z(n1293) );
  CENX1 U1837 ( .A(n1674), .B(n157), .Z(n1307) );
  CENX1 U1838 ( .A(n1684), .B(n156), .Z(n1281) );
  CENX1 U1839 ( .A(n1675), .B(b[24]), .Z(n1306) );
  CENX1 U1840 ( .A(n1564), .B(n104), .Z(n1145) );
  CENX1 U1841 ( .A(n1634), .B(n142), .Z(n1411) );
  CENX1 U1842 ( .A(n1634), .B(n151), .Z(n1406) );
  CENX1 U1843 ( .A(n1662), .B(n152), .Z(n1372) );
  CENX1 U1844 ( .A(n1634), .B(n146), .Z(n1409) );
  CENX1 U1845 ( .A(n1634), .B(n148), .Z(n1408) );
  CENX1 U1846 ( .A(n1654), .B(n152), .Z(n1405) );
  CENX1 U1847 ( .A(n104), .B(a[28]), .Z(n110) );
  CENX1 U1848 ( .A(n1667), .B(n136), .Z(n1350) );
  CENX1 U1849 ( .A(n1654), .B(b[31]), .Z(n1392) );
  CENX1 U1850 ( .A(n1561), .B(n109), .Z(n1140) );
  CENX1 U1851 ( .A(n1666), .B(n138), .Z(n1349) );
  CENX1 U1852 ( .A(n1663), .B(n142), .Z(n1378) );
  CENX1 U1853 ( .A(n1647), .B(a[24]), .Z(n100) );
  CENX1 U1854 ( .A(n109), .B(a[30]), .Z(n114) );
  CENX1 U1855 ( .A(n1659), .B(n154), .Z(n1370) );
  CENX1 U1856 ( .A(n1646), .B(n132), .Z(n1176) );
  CENX1 U1857 ( .A(n1646), .B(n136), .Z(n1174) );
  CENX1 U1858 ( .A(n1645), .B(n142), .Z(n1186) );
  CENX1 U1859 ( .A(n1646), .B(n138), .Z(n1173) );
  CENX1 U1860 ( .A(n1696), .B(n146), .Z(n1220) );
  CENX1 U1861 ( .A(n1696), .B(n148), .Z(n1219) );
  CENX1 U1862 ( .A(n1662), .B(n138), .Z(n1380) );
  CENX1 U1863 ( .A(n1657), .B(b[26]), .Z(n1364) );
  CIVX4 U1864 ( .A(a[0]), .Z(n6) );
  CENX1 U1865 ( .A(n1691), .B(n146), .Z(n1241) );
  CENX1 U1866 ( .A(n1691), .B(n148), .Z(n1240) );
  CENX1 U1867 ( .A(n1677), .B(n152), .Z(n1312) );
  CENX1 U1868 ( .A(n1676), .B(n148), .Z(n1315) );
  CENX1 U1869 ( .A(n1674), .B(n154), .Z(n1310) );
  CENX1 U1870 ( .A(n1676), .B(n146), .Z(n1316) );
  CENX1 U1871 ( .A(n1674), .B(n155), .Z(n1309) );
  CENX1 U1872 ( .A(n1677), .B(n151), .Z(n1313) );
  CENX1 U1873 ( .A(n1670), .B(n146), .Z(n1345) );
  CENX1 U1874 ( .A(n1684), .B(n151), .Z(n1286) );
  CENX1 U1875 ( .A(n1667), .B(n156), .Z(n1337) );
  CENX1 U1876 ( .A(n1684), .B(n146), .Z(n1289) );
  CENX1 U1877 ( .A(n1561), .B(n104), .Z(n1147) );
  CENX1 U1878 ( .A(n1563), .B(n104), .Z(n1146) );
  CENX1 U1879 ( .A(n1562), .B(n104), .Z(n1148) );
  CENX1 U1880 ( .A(n1664), .B(n151), .Z(n1373) );
  CENX1 U1881 ( .A(n1651), .B(n104), .Z(n1149) );
  CENX1 U1882 ( .A(n1667), .B(n157), .Z(n1336) );
  CENX1 U1883 ( .A(n1666), .B(n153), .Z(n1340) );
  CENX1 U1884 ( .A(n1666), .B(b[24]), .Z(n1335) );
  CENX1 U1885 ( .A(n1663), .B(n148), .Z(n1375) );
  CENX1 U1886 ( .A(n1658), .B(b[24]), .Z(n1366) );
  CENX1 U1887 ( .A(n1658), .B(n157), .Z(n1367) );
  CENX1 U1888 ( .A(n1651), .B(n113), .Z(n1137) );
  CENX1 U1889 ( .A(n1666), .B(b[26]), .Z(n1333) );
  CEOX2 U1890 ( .A(n21), .B(a[6]), .Z(n1639) );
  CENX1 U1891 ( .A(n1661), .B(b[29]), .Z(n1361) );
  CNIVX4 U1892 ( .A(n87), .Z(n1646) );
  CEOX1 U1893 ( .A(a[18]), .B(n1645), .Z(n1449) );
  CNIVX4 U1894 ( .A(n93), .Z(n1647) );
  CNIVX4 U1895 ( .A(n99), .Z(n1648) );
  CND2X1 U1896 ( .A(n1444), .B(n110), .Z(n112) );
  CEOXL U1897 ( .A(a[28]), .B(n109), .Z(n1444) );
  CEOX2 U1898 ( .A(n1687), .B(a[12]), .Z(n1623) );
  CEOX1 U1899 ( .A(a[30]), .B(n113), .Z(n1443) );
  CNIVX1 U1900 ( .A(n1056), .Z(n1627) );
  CIVXL U1901 ( .A(n312), .Z(n311) );
  COND2XL U1902 ( .A(n27), .B(n1333), .C(n1332), .D(n24), .Z(n1048) );
  COND2XL U1903 ( .A(n27), .B(n1334), .C(n1333), .D(n24), .Z(n1049) );
  COND2XL U1904 ( .A(n27), .B(n1356), .C(n1355), .D(n24), .Z(n1071) );
  COND2XL U1905 ( .A(n27), .B(n1354), .C(n1353), .D(n24), .Z(n1069) );
  COND2XL U1906 ( .A(n27), .B(n1673), .C(n24), .D(n1360), .Z(n863) );
  COND2XL U1907 ( .A(n1359), .B(n27), .C(n1358), .D(n24), .Z(n1074) );
  COND2XL U1908 ( .A(n27), .B(n1350), .C(n1349), .D(n24), .Z(n1065) );
  COND2XL U1909 ( .A(n27), .B(n1347), .C(n1346), .D(n24), .Z(n1062) );
  COND2XL U1910 ( .A(n27), .B(n1341), .C(n1340), .D(n24), .Z(n1056) );
  COND2XL U1911 ( .A(n27), .B(n1358), .C(n1357), .D(n24), .Z(n1073) );
  COND2XL U1912 ( .A(n27), .B(n1336), .C(n1335), .D(n24), .Z(n1051) );
  COND2XL U1913 ( .A(n27), .B(n1355), .C(n1354), .D(n24), .Z(n1070) );
  CNIVX1 U1914 ( .A(n913), .Z(n1628) );
  CIVX1 U1915 ( .A(n1623), .Z(n1630) );
  CIVX2 U1916 ( .A(n1623), .Z(n1631) );
  CHA1X1 U1917 ( .A(n918), .B(n948), .CO(n668), .S(n669) );
  CIVX2 U1918 ( .A(n1640), .Z(n1675) );
  CFA1XL U1919 ( .A(n897), .B(n977), .CI(n909), .CO(n452), .S(n453) );
  CFA1X1 U1920 ( .A(n854), .B(n1006), .CI(n946), .CO(n626), .S(n627) );
  CIVXL U1921 ( .A(n951), .Z(n1636) );
  CIVX1 U1922 ( .A(n1636), .Z(n1637) );
  CEO3XL U1923 ( .A(n613), .B(n611), .C(n632), .Z(n1638) );
  CIVX1 U1924 ( .A(n1656), .Z(n1655) );
  CND2XL U1925 ( .A(n390), .B(n240), .Z(n172) );
  CIVX1 U1926 ( .A(n240), .Z(n238) );
  CIVXL U1927 ( .A(n239), .Z(n390) );
  CND2XL U1928 ( .A(n391), .B(n250), .Z(n173) );
  CIVX1 U1929 ( .A(n249), .Z(n391) );
  COND2X1 U1930 ( .A(n69), .B(n1226), .C(n1225), .D(n66), .Z(n946) );
  COND2X1 U1931 ( .A(n69), .B(n1228), .C(n1227), .D(n66), .Z(n948) );
  COND2X1 U1932 ( .A(n69), .B(n1223), .C(n1222), .D(n66), .Z(n943) );
  COND2X1 U1933 ( .A(n69), .B(n1225), .C(n1224), .D(n66), .Z(n945) );
  COND2X1 U1934 ( .A(n69), .B(n1230), .C(n1229), .D(n66), .Z(n950) );
  CNR2X2 U1935 ( .A(n609), .B(n630), .Z(n258) );
  CIVX8 U1936 ( .A(n1656), .Z(n1654) );
  CFA1XL U1937 ( .A(n900), .B(n980), .CI(n926), .CO(n534), .S(n535) );
  CIVX2 U1938 ( .A(n1677), .Z(n1640) );
  CENX1 U1939 ( .A(n1651), .B(n1697), .Z(n1233) );
  CENX1 U1940 ( .A(n1559), .B(n1697), .Z(n1234) );
  CENX1 U1941 ( .A(n1697), .B(n151), .Z(n1217) );
  COND2XL U1942 ( .A(n91), .B(n1173), .C(n1172), .D(n89), .Z(n896) );
  COND2XL U1943 ( .A(n91), .B(n1180), .C(n1179), .D(n89), .Z(n903) );
  CNR2IXL U1944 ( .B(n1559), .A(n89), .Z(n907) );
  CND2IXL U1945 ( .B(n1559), .A(n1645), .Z(n1199) );
  COND2XL U1946 ( .A(n53), .B(n1258), .C(n1257), .D(n1597), .Z(n976) );
  CNR2IXL U1947 ( .B(n1559), .A(n1597), .Z(n997) );
  COND2XL U1948 ( .A(n53), .B(n1260), .C(n1259), .D(n1597), .Z(n978) );
  COND2XL U1949 ( .A(n53), .B(n1261), .C(n1260), .D(n1597), .Z(n979) );
  COND2XL U1950 ( .A(n1278), .B(n53), .C(n1277), .D(n1597), .Z(n996) );
  COND2XL U1951 ( .A(n53), .B(n1269), .C(n1268), .D(n1597), .Z(n987) );
  COND2XL U1952 ( .A(n53), .B(n1271), .C(n1270), .D(n1597), .Z(n989) );
  COND2XL U1953 ( .A(n53), .B(n1266), .C(n1265), .D(n1597), .Z(n984) );
  COND2XL U1954 ( .A(n53), .B(n1276), .C(n1275), .D(n1597), .Z(n994) );
  COND2XL U1955 ( .A(n53), .B(n1259), .C(n1258), .D(n1597), .Z(n977) );
  COND2XL U1956 ( .A(n53), .B(n1262), .C(n1261), .D(n1597), .Z(n980) );
  COND2XL U1957 ( .A(n53), .B(n1263), .C(n1262), .D(n1597), .Z(n981) );
  COND2XL U1958 ( .A(n53), .B(n1270), .C(n1269), .D(n1597), .Z(n988) );
  CND2XL U1959 ( .A(n633), .B(n652), .Z(n1641) );
  CND2X1 U1960 ( .A(n633), .B(n635), .Z(n1642) );
  CND2XL U1961 ( .A(n652), .B(n635), .Z(n1643) );
  CND3XL U1962 ( .A(n1641), .B(n1642), .C(n1643), .Z(n630) );
  CIVX1 U1963 ( .A(n30), .Z(n1680) );
  CENX1 U1964 ( .A(n1660), .B(n1562), .Z(n1388) );
  CIVX1 U1965 ( .A(n1665), .Z(n1660) );
  COND2XL U1966 ( .A(n85), .B(n1186), .C(n1185), .D(n82), .Z(n908) );
  COND2XL U1967 ( .A(n85), .B(n1189), .C(n1188), .D(n82), .Z(n911) );
  CNR2IXL U1968 ( .B(n1558), .A(n82), .Z(n921) );
  COND2XL U1969 ( .A(n85), .B(n1188), .C(n1187), .D(n82), .Z(n910) );
  COND2XL U1970 ( .A(n85), .B(n1194), .C(n1193), .D(n82), .Z(n916) );
  COND2XL U1971 ( .A(n85), .B(n1191), .C(n1190), .D(n82), .Z(n913) );
  COND2XL U1972 ( .A(n85), .B(n1193), .C(n1192), .D(n82), .Z(n915) );
  CND2IXL U1973 ( .B(n1559), .A(n1644), .Z(n1216) );
  COND2XL U1974 ( .A(n27), .B(n1353), .C(n1352), .D(n24), .Z(n1068) );
  COND2XL U1975 ( .A(n9), .B(n1656), .C(n6), .D(n1424), .Z(n865) );
  CND2X1 U1976 ( .A(n1136), .B(n865), .Z(n383) );
  CENX1 U1977 ( .A(n1653), .B(b[24]), .Z(n1399) );
  CENX1 U1978 ( .A(n1653), .B(n157), .Z(n1400) );
  CND2IXL U1979 ( .B(n1559), .A(n1634), .Z(n1424) );
  COND2XL U1980 ( .A(n36), .B(n1324), .C(n1323), .D(n33), .Z(n1040) );
  CIVX1 U1981 ( .A(n1679), .Z(n1674) );
  CEOXL U1982 ( .A(n368), .B(n192), .Z(product[5]) );
  CENXL U1983 ( .A(n1659), .B(n155), .Z(n1369) );
  CENXL U1984 ( .A(n1690), .B(n142), .Z(n1243) );
  CND2X4 U1985 ( .A(n1451), .B(n66), .Z(n69) );
  COND2X1 U1986 ( .A(n69), .B(n1227), .C(n1226), .D(n66), .Z(n947) );
  CNR2X1 U1987 ( .A(n651), .B(n670), .Z(n272) );
  CFA1XL U1988 ( .A(n950), .B(n1088), .CI(n1010), .CO(n700), .S(n701) );
  CNIVX1 U1989 ( .A(n120), .Z(n1652) );
  COND2XL U1990 ( .A(n44), .B(n1297), .C(n1296), .D(n42), .Z(n1014) );
  CENX1 U1991 ( .A(n1693), .B(n1563), .Z(n1230) );
  CIVX1 U1992 ( .A(n1673), .Z(n1672) );
  COND2X1 U1993 ( .A(n36), .B(n1325), .C(n1324), .D(n33), .Z(n1041) );
  CENX1 U1994 ( .A(n1669), .B(n1652), .Z(n1358) );
  COND2XL U1995 ( .A(n27), .B(n1357), .C(n1356), .D(n24), .Z(n1072) );
  CHA1XL U1996 ( .A(n859), .B(n1094), .CO(n788), .S(n789) );
  CENX1 U1997 ( .A(n1670), .B(n142), .Z(n1347) );
  CIVX1 U1998 ( .A(n1673), .Z(n1670) );
  COND2XL U1999 ( .A(n53), .B(n1566), .C(n1597), .D(n1279), .Z(n860) );
  CENX1 U2000 ( .A(n189), .B(n357), .Z(product[8]) );
  CENX1 U2001 ( .A(n1663), .B(n146), .Z(n1376) );
  CIVX1 U2002 ( .A(n1665), .Z(n1663) );
  CFA1X1 U2003 ( .A(n984), .B(n894), .CI(n1632), .CO(n622), .S(n623) );
  COND2XL U2004 ( .A(n18), .B(n1369), .C(n15), .D(n1368), .Z(n1083) );
  CIVX2 U2005 ( .A(n1665), .Z(n1658) );
  COND2XL U2006 ( .A(n69), .B(n1218), .C(n1217), .D(n66), .Z(n938) );
  COND2XL U2007 ( .A(n69), .B(n1219), .C(n1218), .D(n66), .Z(n939) );
  COND2XL U2008 ( .A(n69), .B(n1221), .C(n1220), .D(n66), .Z(n941) );
  COND2XL U2009 ( .A(n61), .B(n1692), .C(n1631), .D(n1256), .Z(n859) );
  CNR2IXL U2010 ( .B(n1559), .A(n66), .Z(n955) );
  COND2XL U2011 ( .A(n69), .B(n1220), .C(n1219), .D(n66), .Z(n940) );
  COND2XL U2012 ( .A(n69), .B(n1232), .C(n1231), .D(n66), .Z(n952) );
  COND2XL U2013 ( .A(n69), .B(n1698), .C(n66), .D(n1235), .Z(n858) );
  COND2XL U2014 ( .A(n1234), .B(n69), .C(n1233), .D(n66), .Z(n954) );
  COND2XL U2015 ( .A(n69), .B(n1231), .C(n1230), .D(n66), .Z(n951) );
  CENX1 U2016 ( .A(n1657), .B(b[27]), .Z(n1363) );
  CND2IXL U2017 ( .B(n1559), .A(n1657), .Z(n1391) );
  CIVX2 U2018 ( .A(n1680), .Z(n1676) );
  CNR2X1 U2019 ( .A(n245), .B(n261), .Z(n243) );
  COND1X1 U2020 ( .A(n262), .B(n245), .C(n246), .Z(n244) );
  CND2IXL U2021 ( .B(n1559), .A(n1676), .Z(n1331) );
  CIVX2 U2022 ( .A(n1686), .Z(n1684) );
  CEOXL U2023 ( .A(n199), .B(n166), .Z(product[31]) );
  CND2IXL U2024 ( .B(n1559), .A(n1684), .Z(n1304) );
  CIVX1 U2025 ( .A(n1673), .Z(n1667) );
  CIVX2 U2026 ( .A(n1698), .Z(n1694) );
  CENX1 U2027 ( .A(n1684), .B(n142), .Z(n1291) );
  COND1X1 U2028 ( .A(n226), .B(n1571), .C(n219), .Z(n217) );
  CIVX1 U2029 ( .A(n1673), .Z(n1666) );
  COND2XL U2030 ( .A(n18), .B(n1362), .C(n15), .D(n1361), .Z(n1076) );
  COND2XL U2031 ( .A(n18), .B(n1387), .C(n15), .D(n1386), .Z(n1101) );
  COND2XL U2032 ( .A(n18), .B(n1363), .C(n15), .D(n1362), .Z(n1077) );
  COND2XL U2033 ( .A(n18), .B(n1385), .C(n15), .D(n1384), .Z(n1099) );
  COND2XL U2034 ( .A(n1390), .B(n18), .C(n15), .D(n1389), .Z(n1104) );
  COND2XL U2035 ( .A(n18), .B(n1388), .C(n15), .D(n1387), .Z(n1102) );
  COND2XL U2036 ( .A(n18), .B(n1383), .C(n15), .D(n1382), .Z(n1097) );
  COND2XL U2037 ( .A(n18), .B(n1386), .C(n15), .D(n1385), .Z(n1100) );
  COND2XL U2038 ( .A(n18), .B(n1365), .C(n15), .D(n1364), .Z(n1079) );
  COND2XL U2039 ( .A(n18), .B(n1665), .C(n15), .D(n1391), .Z(n864) );
  COND2XL U2040 ( .A(n18), .B(n1364), .C(n15), .D(n1363), .Z(n1078) );
  COND2XL U2041 ( .A(n18), .B(n1382), .C(n15), .D(n1381), .Z(n1096) );
  COND2XL U2042 ( .A(n18), .B(n1384), .C(n15), .D(n1383), .Z(n1098) );
  COND2XL U2043 ( .A(n18), .B(n1379), .C(n15), .D(n1378), .Z(n1093) );
  COND2XL U2044 ( .A(n18), .B(n1381), .C(n15), .D(n1380), .Z(n1095) );
  COND2XL U2045 ( .A(n18), .B(n1376), .C(n15), .D(n1375), .Z(n1090) );
  COND2XL U2046 ( .A(n18), .B(n1367), .C(n15), .D(n1366), .Z(n1081) );
  COND2XL U2047 ( .A(n18), .B(n1380), .C(n15), .D(n1379), .Z(n1094) );
  COND2XL U2048 ( .A(n18), .B(n1370), .C(n15), .D(n1369), .Z(n1084) );
  CIVXL U2049 ( .A(n1572), .Z(n387) );
  CNR2X1 U2050 ( .A(n218), .B(n223), .Z(n216) );
  COAN1X1 U2051 ( .A(n259), .B(n249), .C(n250), .Z(n246) );
  CIVX2 U2052 ( .A(n1665), .Z(n1664) );
  CENX1 U2053 ( .A(n1676), .B(n138), .Z(n1320) );
  CND2X1 U2054 ( .A(n391), .B(n392), .Z(n245) );
  CIVX2 U2055 ( .A(n1698), .Z(n1697) );
  CIVX4 U2056 ( .A(n12), .Z(n1665) );
  CANR1X2 U2057 ( .A(n243), .B(n279), .C(n244), .Z(n242) );
  CND2X4 U2058 ( .A(n1458), .B(n6), .Z(n9) );
  CENX4 U2059 ( .A(n1654), .B(a[2]), .Z(n15) );
  CND2X4 U2060 ( .A(n1457), .B(n15), .Z(n18) );
  CND2X4 U2061 ( .A(n1456), .B(n24), .Z(n27) );
  CND2X4 U2062 ( .A(n1455), .B(n33), .Z(n36) );
  CND2X4 U2063 ( .A(n1452), .B(n1629), .Z(n61) );
  CENX4 U2064 ( .A(n1690), .B(a[14]), .Z(n66) );
  CIVXL U2065 ( .A(n1665), .Z(n1657) );
  CIVXL U2066 ( .A(n1665), .Z(n1659) );
  CIVXL U2067 ( .A(n1665), .Z(n1662) );
  CIVXL U2068 ( .A(n1673), .Z(n1668) );
  CIVXL U2069 ( .A(n1673), .Z(n1669) );
  CIVXL U2070 ( .A(n1673), .Z(n1671) );
  CIVXL U2071 ( .A(n30), .Z(n1678) );
  CIVXL U2072 ( .A(n1685), .Z(n1681) );
  CIVXL U2073 ( .A(n1685), .Z(n1683) );
  CIVXL U2074 ( .A(n1698), .Z(n1696) );
  CIVX2 U2075 ( .A(n374), .Z(n412) );
  CIVX2 U2076 ( .A(n358), .Z(n408) );
  CIVX2 U2077 ( .A(n336), .Z(n404) );
  CIVX2 U2078 ( .A(n333), .Z(n403) );
  CIVX2 U2079 ( .A(n322), .Z(n401) );
  CIVX2 U2080 ( .A(n295), .Z(n397) );
  CIVX2 U2081 ( .A(n234), .Z(n389) );
  CIVX2 U2082 ( .A(n223), .Z(n388) );
  CIVX2 U2083 ( .A(n383), .Z(n381) );
  CIVX2 U2084 ( .A(n380), .Z(n378) );
  CIVX2 U2085 ( .A(n372), .Z(n370) );
  CIVX2 U2086 ( .A(n364), .Z(n362) );
  CIVX2 U2087 ( .A(n356), .Z(n354) );
  CIVX2 U2088 ( .A(n352), .Z(n351) );
  CIVX2 U2089 ( .A(n350), .Z(n348) );
  CIVX2 U2090 ( .A(n345), .Z(n343) );
  CIVX2 U2091 ( .A(n339), .Z(n338) );
  CIVX2 U2092 ( .A(n328), .Z(n326) );
  CIVX2 U2093 ( .A(n327), .Z(n402) );
  CIVX2 U2094 ( .A(n318), .Z(n316) );
  CIVX2 U2095 ( .A(n305), .Z(n399) );
  CIVX2 U2096 ( .A(n303), .Z(n301) );
  CIVX2 U2097 ( .A(n290), .Z(n288) );
  CIVX2 U2098 ( .A(n285), .Z(n283) );
  CIVX2 U2099 ( .A(n272), .Z(n394) );
  CIVX2 U2100 ( .A(n270), .Z(n268) );
  CIVX2 U2101 ( .A(n261), .Z(n263) );
  CIVX2 U2102 ( .A(n259), .Z(n257) );
  CIVX2 U2103 ( .A(n258), .Z(n392) );
  CIVX2 U2104 ( .A(n242), .Z(n241) );
  CIVX2 U2105 ( .A(n229), .Z(n231) );
  CIVX2 U2106 ( .A(n212), .Z(n210) );
  CIVX2 U2107 ( .A(n207), .Z(n205) );
  CIVX2 U2108 ( .A(n206), .Z(n385) );
  CIVX2 U2109 ( .A(n1647), .Z(n1472) );
  CIVX2 U2110 ( .A(n1648), .Z(n1471) );
  CIVX2 U2111 ( .A(n104), .Z(n1470) );
  CIVX2 U2112 ( .A(n109), .Z(n1469) );
  CIVX2 U2113 ( .A(n113), .Z(n1468) );
endmodule


module calc_DW_mult_uns_16 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n3, n6, n9, n12, n15, n18, n21, n24, n27, n30, n33, n36, n39, n42,
         n44, n48, n50, n53, n55, n58, n61, n63, n66, n69, n71, n74, n77, n79,
         n82, n85, n87, n89, n91, n93, n95, n97, n99, n100, n102, n104, n105,
         n107, n109, n110, n112, n113, n114, n115, n116, n120, n122, n124,
         n126, n128, n130, n132, n134, n136, n138, n140, n142, n144, n146,
         n148, n150, n151, n152, n153, n154, n155, n156, n157, n169, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n198, n199, n205, n207, n208, n210, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n226, n227, n228,
         n229, n234, n235, n236, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n248, n250, n251, n252, n253, n257, n259, n260, n261,
         n262, n263, n264, n268, n270, n271, n272, n273, n275, n278, n279,
         n280, n281, n283, n285, n286, n288, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n301, n303, n304, n305, n306, n308,
         n312, n313, n314, n316, n318, n319, n320, n321, n322, n323, n324,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n343, n345, n346, n348, n350, n351,
         n352, n354, n356, n357, n358, n359, n360, n362, n364, n365, n366,
         n367, n368, n370, n372, n373, n374, n375, n376, n378, n380, n381,
         n383, n388, n389, n390, n394, n397, n399, n401, n402, n403, n404,
         n412, n415, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1455, n1457,
         n1458, n1468, n1469, n1470, n1471, n1475, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724;
  assign n3 = a[1];
  assign n12 = a[3];
  assign n21 = a[5];
  assign n30 = a[7];
  assign n39 = a[9];
  assign n48 = a[11];
  assign n55 = a[13];
  assign n63 = a[15];
  assign n71 = a[17];
  assign n79 = a[19];
  assign n87 = a[21];
  assign n93 = a[23];
  assign n99 = a[25];
  assign n104 = a[27];
  assign n109 = a[29];
  assign n113 = a[31];
  assign n116 = b[0];
  assign n120 = b[1];
  assign n122 = b[2];
  assign n124 = b[3];
  assign n126 = b[4];
  assign n128 = b[5];
  assign n130 = b[6];
  assign n132 = b[7];
  assign n134 = b[8];
  assign n136 = b[9];
  assign n138 = b[10];
  assign n140 = b[11];
  assign n142 = b[12];
  assign n144 = b[13];
  assign n146 = b[14];
  assign n148 = b[15];
  assign n150 = b[16];
  assign n151 = b[17];
  assign n152 = b[18];
  assign n153 = b[19];
  assign n154 = b[20];
  assign n155 = b[21];
  assign n156 = b[22];
  assign n157 = b[23];

  CEO3X2 U410 ( .A(n420), .B(n438), .C(n419), .Z(n417) );
  CEO3X2 U411 ( .A(n422), .B(n421), .C(n440), .Z(n418) );
  CEO3X2 U412 ( .A(n444), .B(n423), .C(n442), .Z(n419) );
  CEO3X2 U413 ( .A(n425), .B(n424), .C(n446), .Z(n420) );
  CEO3X2 U416 ( .A(n456), .B(n429), .C(n454), .Z(n423) );
  CEO3X2 U417 ( .A(n998), .B(n1106), .C(n1076), .Z(n424) );
  CEO3X2 U418 ( .A(n956), .B(n1048), .C(n866), .Z(n425) );
  CEO3X2 U419 ( .A(n908), .B(n938), .C(n1022), .Z(n426) );
  CEO3X2 U421 ( .A(n878), .B(n868), .C(n850), .Z(n428) );
  CFA1X1 U423 ( .A(n435), .B(n433), .CI(n460), .CO(n430), .S(n431) );
  CFA1X1 U424 ( .A(n439), .B(n462), .CI(n437), .CO(n432), .S(n433) );
  CFA1X1 U425 ( .A(n441), .B(n464), .CI(n466), .CO(n434), .S(n435) );
  CFA1X1 U426 ( .A(n445), .B(n443), .CI(n468), .CO(n436), .S(n437) );
  CFA1X1 U427 ( .A(n472), .B(n447), .CI(n470), .CO(n438), .S(n439) );
  CFA1X1 U428 ( .A(n451), .B(n449), .CI(n474), .CO(n440), .S(n441) );
  CFA1X1 U429 ( .A(n457), .B(n453), .CI(n455), .CO(n442), .S(n443) );
  CFA1X1 U430 ( .A(n480), .B(n476), .CI(n478), .CO(n444), .S(n445) );
  CFA1X1 U431 ( .A(n1023), .B(n482), .CI(n484), .CO(n446), .S(n447) );
  CFA1X1 U432 ( .A(n957), .B(n1049), .CI(n1107), .CO(n448), .S(n449) );
  CFA1X1 U433 ( .A(n939), .B(n1077), .CI(n999), .CO(n450), .S(n451) );
  CFA1X1 U434 ( .A(n897), .B(n977), .CI(n909), .CO(n452), .S(n453) );
  CFA1X1 U435 ( .A(n869), .B(n923), .CI(n887), .CO(n454), .S(n455) );
  CFA1X1 U436 ( .A(n867), .B(n879), .CI(n873), .CO(n456), .S(n457) );
  CFA1X1 U437 ( .A(n463), .B(n461), .CI(n488), .CO(n458), .S(n459) );
  CFA1X1 U438 ( .A(n467), .B(n490), .CI(n465), .CO(n460), .S(n461) );
  CFA1X1 U439 ( .A(n469), .B(n492), .CI(n494), .CO(n462), .S(n463) );
  CFA1X1 U440 ( .A(n473), .B(n471), .CI(n496), .CO(n464), .S(n465) );
  CFA1X1 U441 ( .A(n475), .B(n498), .CI(n500), .CO(n466), .S(n467) );
  CFA1X1 U442 ( .A(n481), .B(n477), .CI(n479), .CO(n468), .S(n469) );
  CFA1X1 U443 ( .A(n502), .B(n483), .CI(n504), .CO(n470), .S(n471) );
  CFA1X1 U444 ( .A(n510), .B(n506), .CI(n508), .CO(n472), .S(n473) );
  CFA1X1 U445 ( .A(n1024), .B(n485), .CI(n1108), .CO(n474), .S(n475) );
  CFA1X1 U447 ( .A(n940), .B(n870), .CI(n1561), .CO(n478), .S(n479) );
  CFA1X1 U448 ( .A(n851), .B(n978), .CI(n924), .CO(n480), .S(n481) );
  CFA1X1 U449 ( .A(n874), .B(n910), .CI(n898), .CO(n482), .S(n483) );
  CHA1X1 U450 ( .A(n880), .B(n888), .CO(n484), .S(n485) );
  CFA1X1 U452 ( .A(n495), .B(n516), .CI(n493), .CO(n488), .S(n489) );
  CFA1X1 U453 ( .A(n497), .B(n518), .CI(n520), .CO(n490), .S(n491) );
  CFA1X1 U454 ( .A(n501), .B(n499), .CI(n522), .CO(n492), .S(n493) );
  CFA1X1 U455 ( .A(n503), .B(n524), .CI(n526), .CO(n494), .S(n495) );
  CFA1X1 U456 ( .A(n509), .B(n505), .CI(n507), .CO(n496), .S(n497) );
  CFA1X1 U457 ( .A(n530), .B(n511), .CI(n528), .CO(n498), .S(n499) );
  CFA1X1 U458 ( .A(n536), .B(n534), .CI(n532), .CO(n500), .S(n501) );
  CFA1X1 U459 ( .A(n979), .B(n1109), .CI(n1001), .CO(n502), .S(n503) );
  CFA1X1 U461 ( .A(n911), .B(n1025), .CI(n925), .CO(n506), .S(n507) );
  CFA1X1 U462 ( .A(n889), .B(n941), .CI(n899), .CO(n508), .S(n509) );
  CFA1X1 U463 ( .A(n871), .B(n875), .CI(n881), .CO(n510), .S(n511) );
  CFA1X1 U464 ( .A(n517), .B(n515), .CI(n540), .CO(n512), .S(n513) );
  CFA1X1 U465 ( .A(n521), .B(n542), .CI(n519), .CO(n514), .S(n515) );
  CFA1X1 U466 ( .A(n546), .B(n544), .CI(n523), .CO(n516), .S(n517) );
  CFA1X1 U467 ( .A(n527), .B(n525), .CI(n548), .CO(n518), .S(n519) );
  CFA1X1 U468 ( .A(n535), .B(n550), .CI(n529), .CO(n520), .S(n521) );
  CFA1X1 U469 ( .A(n552), .B(n531), .CI(n533), .CO(n522), .S(n523) );
  CFA1X1 U470 ( .A(n558), .B(n554), .CI(n556), .CO(n524), .S(n525) );
  CFA1X1 U471 ( .A(n1110), .B(n560), .CI(n537), .CO(n526), .S(n527) );
  CFA1X1 U473 ( .A(n942), .B(n876), .CI(n1002), .CO(n530), .S(n531) );
  CFA1X1 U474 ( .A(n852), .B(n960), .CI(n912), .CO(n532), .S(n533) );
  CFA1X1 U475 ( .A(n900), .B(n980), .CI(n926), .CO(n534), .S(n535) );
  CFA1X1 U477 ( .A(n543), .B(n541), .CI(n564), .CO(n538), .S(n539) );
  CFA1X1 U478 ( .A(n568), .B(n566), .CI(n545), .CO(n540), .S(n541) );
  CFA1X1 U479 ( .A(n570), .B(n547), .CI(n549), .CO(n542), .S(n543) );
  CFA1X1 U480 ( .A(n574), .B(n551), .CI(n572), .CO(n544), .S(n545) );
  CFA1X1 U481 ( .A(n557), .B(n553), .CI(n555), .CO(n546), .S(n547) );
  CFA1X1 U482 ( .A(n578), .B(n559), .CI(n561), .CO(n548), .S(n549) );
  CFA1X1 U483 ( .A(n582), .B(n576), .CI(n580), .CO(n550), .S(n551) );
  CFA1X1 U484 ( .A(n1003), .B(n584), .CI(n1111), .CO(n552), .S(n553) );
  CFA1X1 U485 ( .A(n961), .B(n1081), .CI(n1053), .CO(n554), .S(n555) );
  CFA1X1 U486 ( .A(n913), .B(n1027), .CI(n943), .CO(n556), .S(n557) );
  CFA1X1 U487 ( .A(n901), .B(n981), .CI(n927), .CO(n558), .S(n559) );
  CFA1X1 U488 ( .A(n877), .B(n1617), .CI(n883), .CO(n560), .S(n561) );
  CFA1X1 U489 ( .A(n567), .B(n565), .CI(n588), .CO(n562), .S(n563) );
  CFA1X1 U490 ( .A(n592), .B(n590), .CI(n569), .CO(n564), .S(n565) );
  CFA1X1 U491 ( .A(n594), .B(n571), .CI(n573), .CO(n566), .S(n567) );
  CFA1X1 U492 ( .A(n598), .B(n575), .CI(n596), .CO(n568), .S(n569) );
  CFA1X1 U493 ( .A(n581), .B(n577), .CI(n579), .CO(n570), .S(n571) );
  CFA1X1 U495 ( .A(n585), .B(n604), .CI(n606), .CO(n574), .S(n575) );
  CFA1X1 U496 ( .A(n1004), .B(n1082), .CI(n1112), .CO(n576), .S(n577) );
  CFA1X1 U497 ( .A(n962), .B(n884), .CI(n1054), .CO(n578), .S(n579) );
  CFA1X1 U498 ( .A(n914), .B(n1028), .CI(n944), .CO(n580), .S(n581) );
  CFA1X1 U499 ( .A(n902), .B(n982), .CI(n928), .CO(n582), .S(n583) );
  CHA1X1 U500 ( .A(n892), .B(n853), .CO(n584), .S(n585) );
  CFA1X1 U501 ( .A(n591), .B(n589), .CI(n610), .CO(n586), .S(n587) );
  CFA1X1 U502 ( .A(n614), .B(n593), .CI(n612), .CO(n588), .S(n589) );
  CFA1X1 U503 ( .A(n616), .B(n595), .CI(n597), .CO(n590), .S(n591) );
  CFA1X1 U504 ( .A(n620), .B(n599), .CI(n618), .CO(n592), .S(n593) );
  CFA1X1 U505 ( .A(n605), .B(n601), .CI(n603), .CO(n594), .S(n595) );
  CFA1X1 U506 ( .A(n624), .B(n607), .CI(n622), .CO(n596), .S(n597) );
  CFA1X1 U507 ( .A(n1005), .B(n626), .CI(n628), .CO(n598), .S(n599) );
  CFA1X1 U508 ( .A(n983), .B(n1113), .CI(n1055), .CO(n600), .S(n601) );
  CFA1X1 U509 ( .A(n929), .B(n1083), .CI(n963), .CO(n602), .S(n603) );
  CFA1X1 U510 ( .A(n1615), .B(n1029), .CI(n945), .CO(n604), .S(n605) );
  CFA1X1 U511 ( .A(n885), .B(n903), .CI(n893), .CO(n606), .S(n607) );
  CFA1X1 U512 ( .A(n613), .B(n611), .CI(n632), .CO(n608), .S(n609) );
  CFA1X1 U513 ( .A(n617), .B(n634), .CI(n615), .CO(n610), .S(n611) );
  CFA1X1 U515 ( .A(n623), .B(n640), .CI(n621), .CO(n614), .S(n615) );
  CFA1X1 U516 ( .A(n642), .B(n625), .CI(n627), .CO(n616), .S(n617) );
  CFA1X1 U517 ( .A(n648), .B(n646), .CI(n644), .CO(n618), .S(n619) );
  CFA1X1 U518 ( .A(n1114), .B(n629), .CI(n1573), .CO(n620), .S(n621) );
  CFA1X1 U519 ( .A(n984), .B(n894), .CI(n1084), .CO(n622), .S(n623) );
  CFA1X1 U521 ( .A(n854), .B(n1006), .CI(n946), .CO(n626), .S(n627) );
  CHA1X1 U522 ( .A(n904), .B(n930), .CO(n628), .S(n629) );
  CFA1X1 U524 ( .A(n639), .B(n654), .CI(n637), .CO(n632), .S(n633) );
  CFA1X1 U525 ( .A(n658), .B(n656), .CI(n641), .CO(n634), .S(n635) );
  CFA1X1 U526 ( .A(n645), .B(n660), .CI(n643), .CO(n636), .S(n637) );
  CFA1X1 U528 ( .A(n668), .B(n664), .CI(n666), .CO(n640), .S(n641) );
  CFA1X1 U529 ( .A(n985), .B(n1115), .CI(n1031), .CO(n642), .S(n643) );
  CFA1X1 U530 ( .A(n947), .B(n1057), .CI(n1007), .CO(n644), .S(n645) );
  CFA1X1 U531 ( .A(n931), .B(n1085), .CI(n965), .CO(n646), .S(n647) );
  CFA1X1 U532 ( .A(n895), .B(n1611), .CI(n905), .CO(n648), .S(n649) );
  CFA1X1 U533 ( .A(n655), .B(n653), .CI(n672), .CO(n650), .S(n651) );
  CFA1X1 U534 ( .A(n659), .B(n674), .CI(n657), .CO(n652), .S(n653) );
  CFA1X1 U535 ( .A(n678), .B(n676), .CI(n661), .CO(n654), .S(n655) );
  CFA1X1 U536 ( .A(n665), .B(n663), .CI(n680), .CO(n656), .S(n657) );
  CFA1X1 U537 ( .A(n684), .B(n667), .CI(n682), .CO(n658), .S(n659) );
  CFA1X1 U538 ( .A(n1032), .B(n669), .CI(n686), .CO(n660), .S(n661) );
  CFA1X1 U539 ( .A(n1008), .B(n1116), .CI(n1058), .CO(n662), .S(n663) );
  CFA1X1 U540 ( .A(n855), .B(n1086), .CI(n986), .CO(n664), .S(n665) );
  CFA1X1 U541 ( .A(n932), .B(n906), .CI(n966), .CO(n666), .S(n667) );
  CHA1X1 U542 ( .A(n948), .B(n918), .CO(n668), .S(n669) );
  CFA1X1 U543 ( .A(n675), .B(n673), .CI(n690), .CO(n670), .S(n671) );
  CFA1X1 U544 ( .A(n679), .B(n692), .CI(n677), .CO(n672), .S(n673) );
  CFA1X1 U545 ( .A(n681), .B(n694), .CI(n696), .CO(n674), .S(n675) );
  CFA1X1 U546 ( .A(n687), .B(n683), .CI(n685), .CO(n676), .S(n677) );
  CFA1X1 U547 ( .A(n702), .B(n698), .CI(n700), .CO(n678), .S(n679) );
  CFA1X1 U548 ( .A(n987), .B(n704), .CI(n1033), .CO(n680), .S(n681) );
  CFA1X1 U549 ( .A(n967), .B(n1059), .CI(n1117), .CO(n682), .S(n683) );
  CFA1X1 U551 ( .A(n907), .B(n933), .CI(n919), .CO(n686), .S(n687) );
  CFA1X1 U552 ( .A(n693), .B(n691), .CI(n708), .CO(n688), .S(n689) );
  CFA1X1 U553 ( .A(n697), .B(n710), .CI(n695), .CO(n690), .S(n691) );
  CFA1X1 U554 ( .A(n699), .B(n712), .CI(n714), .CO(n692), .S(n693) );
  CFA1X1 U555 ( .A(n718), .B(n701), .CI(n703), .CO(n694), .S(n695) );
  CFA1X1 U556 ( .A(n705), .B(n716), .CI(n720), .CO(n696), .S(n697) );
  CFA1X1 U557 ( .A(n1034), .B(n1118), .CI(n1060), .CO(n698), .S(n699) );
  CFA1X1 U558 ( .A(n950), .B(n1088), .CI(n1010), .CO(n700), .S(n701) );
  CFA1X1 U559 ( .A(n856), .B(n1613), .CI(n968), .CO(n702), .S(n703) );
  CHA1X1 U560 ( .A(n934), .B(n988), .CO(n704), .S(n705) );
  CFA1X1 U561 ( .A(n711), .B(n709), .CI(n724), .CO(n706), .S(n707) );
  CFA1X1 U562 ( .A(n715), .B(n726), .CI(n713), .CO(n708), .S(n709) );
  CFA1X1 U563 ( .A(n717), .B(n728), .CI(n730), .CO(n710), .S(n711) );
  CFA1X1 U564 ( .A(n732), .B(n719), .CI(n721), .CO(n712), .S(n713) );
  CFA1X1 U565 ( .A(n1011), .B(n734), .CI(n736), .CO(n714), .S(n715) );
  CFA1X1 U566 ( .A(n989), .B(n1119), .CI(n1035), .CO(n716), .S(n717) );
  CFA1X1 U567 ( .A(n969), .B(n1089), .CI(n1061), .CO(n718), .S(n719) );
  CFA1X1 U568 ( .A(n921), .B(n951), .CI(n935), .CO(n720), .S(n721) );
  CFA1X1 U569 ( .A(n727), .B(n725), .CI(n740), .CO(n722), .S(n723) );
  CFA1X1 U570 ( .A(n744), .B(n742), .CI(n729), .CO(n724), .S(n725) );
  CFA1X1 U571 ( .A(n735), .B(n731), .CI(n733), .CO(n726), .S(n727) );
  CFA1X1 U572 ( .A(n750), .B(n748), .CI(n746), .CO(n728), .S(n729) );
  CFA1X1 U574 ( .A(n970), .B(n1090), .CI(n1120), .CO(n732), .S(n733) );
  CFA1X1 U575 ( .A(n952), .B(n936), .CI(n990), .CO(n734), .S(n735) );
  CHA1X1 U576 ( .A(n857), .B(n1012), .CO(n736), .S(n737) );
  CFA1X1 U577 ( .A(n743), .B(n741), .CI(n754), .CO(n738), .S(n739) );
  CFA1X1 U578 ( .A(n758), .B(n756), .CI(n745), .CO(n740), .S(n741) );
  CFA1X1 U579 ( .A(n751), .B(n747), .CI(n749), .CO(n742), .S(n743) );
  CFA1X1 U580 ( .A(n764), .B(n760), .CI(n762), .CO(n744), .S(n745) );
  CFA1X1 U582 ( .A(n991), .B(n1091), .CI(n1063), .CO(n748), .S(n749) );
  CFA1X1 U583 ( .A(n937), .B(n971), .CI(n953), .CO(n750), .S(n751) );
  CFA1X1 U584 ( .A(n757), .B(n755), .CI(n768), .CO(n752), .S(n753) );
  CFA1X1 U585 ( .A(n772), .B(n759), .CI(n770), .CO(n754), .S(n755) );
  CFA1X1 U586 ( .A(n774), .B(n761), .CI(n763), .CO(n756), .S(n757) );
  CFA1X1 U587 ( .A(n1038), .B(n776), .CI(n765), .CO(n758), .S(n759) );
  CFA1X1 U588 ( .A(n992), .B(n1092), .CI(n1064), .CO(n760), .S(n761) );
  CFA1X1 U589 ( .A(n972), .B(n954), .CI(n1122), .CO(n762), .S(n763) );
  CHA1X1 U590 ( .A(n858), .B(n1014), .CO(n764), .S(n765) );
  CFA1X1 U591 ( .A(n771), .B(n769), .CI(n780), .CO(n766), .S(n767) );
  CFA1X1 U592 ( .A(n775), .B(n782), .CI(n773), .CO(n768), .S(n769) );
  CFA1X1 U593 ( .A(n784), .B(n777), .CI(n786), .CO(n770), .S(n771) );
  CFA1X1 U595 ( .A(n1015), .B(n1093), .CI(n1123), .CO(n774), .S(n775) );
  CFA1X1 U596 ( .A(n955), .B(n993), .CI(n973), .CO(n776), .S(n777) );
  CFA1X1 U597 ( .A(n783), .B(n781), .CI(n792), .CO(n778), .S(n779) );
  CFA1X1 U598 ( .A(n787), .B(n794), .CI(n785), .CO(n780), .S(n781) );
  CFA1X1 U599 ( .A(n789), .B(n796), .CI(n798), .CO(n782), .S(n783) );
  CFA1X1 U600 ( .A(n1016), .B(n1066), .CI(n1040), .CO(n784), .S(n785) );
  CFA1X1 U601 ( .A(n994), .B(n974), .CI(n1124), .CO(n786), .S(n787) );
  CHA1X1 U602 ( .A(n859), .B(n1094), .CO(n788), .S(n789) );
  CFA1X1 U603 ( .A(n802), .B(n793), .CI(n795), .CO(n790), .S(n791) );
  CFA1X1 U604 ( .A(n799), .B(n804), .CI(n797), .CO(n792), .S(n793) );
  CFA1X1 U605 ( .A(n1125), .B(n806), .CI(n808), .CO(n794), .S(n795) );
  CFA1X1 U606 ( .A(n1041), .B(n1095), .CI(n1067), .CO(n796), .S(n797) );
  CFA1X1 U607 ( .A(n975), .B(n1017), .CI(n995), .CO(n798), .S(n799) );
  CFA1X1 U608 ( .A(n805), .B(n803), .CI(n812), .CO(n800), .S(n801) );
  CFA1X1 U609 ( .A(n816), .B(n807), .CI(n814), .CO(n802), .S(n803) );
  CFA1X1 U610 ( .A(n1042), .B(n809), .CI(n1068), .CO(n804), .S(n805) );
  CFA1X1 U611 ( .A(n1557), .B(n1096), .CI(n1126), .CO(n806), .S(n807) );
  CFA1X1 U613 ( .A(n815), .B(n813), .CI(n820), .CO(n810), .S(n811) );
  CFA1X1 U614 ( .A(n824), .B(n817), .CI(n822), .CO(n812), .S(n813) );
  CFA1X1 U615 ( .A(n1127), .B(n1097), .CI(n1069), .CO(n814), .S(n815) );
  CFA1X1 U616 ( .A(n997), .B(n1043), .CI(n1019), .CO(n816), .S(n817) );
  CFA1X1 U617 ( .A(n828), .B(n821), .CI(n823), .CO(n818), .S(n819) );
  CFA1X1 U618 ( .A(n1128), .B(n830), .CI(n825), .CO(n820), .S(n821) );
  CFA1X1 U619 ( .A(n1044), .B(n1098), .CI(n1070), .CO(n822), .S(n823) );
  CHA1X1 U620 ( .A(n861), .B(n1020), .CO(n824), .S(n825) );
  CFA1X1 U621 ( .A(n834), .B(n829), .CI(n831), .CO(n826), .S(n827) );
  CFA1X1 U622 ( .A(n1071), .B(n836), .CI(n1099), .CO(n828), .S(n829) );
  CFA1X1 U624 ( .A(n837), .B(n835), .CI(n840), .CO(n832), .S(n833) );
  CHA1X1 U626 ( .A(n862), .B(n1046), .CO(n836), .S(n837) );
  CFA1X1 U627 ( .A(n1101), .B(n841), .CI(n844), .CO(n838), .S(n839) );
  CFA1X1 U628 ( .A(n1047), .B(n1073), .CI(n1131), .CO(n840), .S(n841) );
  CFA1X1 U629 ( .A(n1132), .B(n845), .CI(n1102), .CO(n842), .S(n843) );
  CHA1X1 U630 ( .A(n863), .B(n1074), .CO(n844), .S(n845) );
  CFA1X1 U631 ( .A(n1075), .B(n1103), .CI(n1133), .CO(n846), .S(n847) );
  CHA1X1 U632 ( .A(n1134), .B(n864), .CO(n848), .S(n849) );
  COND2X1 U633 ( .A(n1139), .B(n114), .C(n1468), .D(n115), .Z(n850) );
  COND2X1 U634 ( .A(n1138), .B(n115), .C(n114), .D(n1137), .Z(n866) );
  CND2IX1 U638 ( .B(n1687), .A(n113), .Z(n1139) );
  COND2X1 U639 ( .A(n1144), .B(n110), .C(n1469), .D(n112), .Z(n851) );
  COND2X1 U640 ( .A(n112), .B(n1141), .C(n110), .D(n1140), .Z(n868) );
  COND2X1 U641 ( .A(n112), .B(n1142), .C(n110), .D(n1141), .Z(n869) );
  COND2X1 U642 ( .A(n1143), .B(n112), .C(n110), .D(n1142), .Z(n870) );
  COND2X1 U650 ( .A(n107), .B(n1146), .C(n105), .D(n1145), .Z(n872) );
  COND2X1 U651 ( .A(n107), .B(n1147), .C(n105), .D(n1146), .Z(n873) );
  COND2X1 U652 ( .A(n107), .B(n1148), .C(n105), .D(n1147), .Z(n874) );
  COND2X1 U653 ( .A(n1149), .B(n107), .C(n105), .D(n1148), .Z(n875) );
  COND2X1 U654 ( .A(n1150), .B(n107), .C(n105), .D(n1149), .Z(n876) );
  CND2IX1 U662 ( .B(n1687), .A(n104), .Z(n1151) );
  COND2X1 U664 ( .A(n102), .B(n1153), .C(n1609), .D(n1152), .Z(n878) );
  COND2X1 U665 ( .A(n102), .B(n1154), .C(n1609), .D(n1153), .Z(n879) );
  COND2X1 U667 ( .A(n102), .B(n1156), .C(n1609), .D(n1155), .Z(n881) );
  COND2X1 U669 ( .A(n102), .B(n1158), .C(n1609), .D(n1157), .Z(n883) );
  COND2X1 U670 ( .A(n1159), .B(n102), .C(n1609), .D(n1158), .Z(n884) );
  CND2IX1 U680 ( .B(n1687), .A(n1685), .Z(n1160) );
  COND2X1 U683 ( .A(n97), .B(n1163), .C(n1162), .D(n95), .Z(n887) );
  COND2X1 U685 ( .A(n97), .B(n1165), .C(n1164), .D(n95), .Z(n889) );
  CND2IX1 U702 ( .B(n1687), .A(n1684), .Z(n1171) );
  COND2X1 U703 ( .A(n1184), .B(n89), .C(n1628), .D(n91), .Z(n855) );
  COND2X1 U704 ( .A(n91), .B(n1173), .C(n1172), .D(n89), .Z(n896) );
  COND2X1 U705 ( .A(n91), .B(n1174), .C(n1173), .D(n89), .Z(n897) );
  COND2X1 U706 ( .A(n91), .B(n1175), .C(n1174), .D(n89), .Z(n898) );
  COND2X1 U707 ( .A(n91), .B(n1176), .C(n1175), .D(n89), .Z(n899) );
  COND2X1 U708 ( .A(n91), .B(n1177), .C(n1176), .D(n89), .Z(n900) );
  COND2X1 U709 ( .A(n91), .B(n1178), .C(n1177), .D(n89), .Z(n901) );
  COND2X1 U710 ( .A(n91), .B(n1179), .C(n1178), .D(n89), .Z(n902) );
  COND2X1 U711 ( .A(n91), .B(n1180), .C(n1179), .D(n89), .Z(n903) );
  COND2X1 U712 ( .A(n91), .B(n1181), .C(n89), .D(n1180), .Z(n904) );
  COND2X1 U713 ( .A(n91), .B(n1182), .C(n89), .D(n1181), .Z(n905) );
  COND2X1 U714 ( .A(n1183), .B(n91), .C(n89), .D(n1182), .Z(n906) );
  COND2X1 U729 ( .A(n85), .B(n1600), .C(n1666), .D(n1199), .Z(n856) );
  COND2X1 U734 ( .A(n85), .B(n1190), .C(n1189), .D(n1666), .Z(n912) );
  COND2X1 U736 ( .A(n85), .B(n1192), .C(n1191), .D(n1666), .Z(n914) );
  COND2X1 U740 ( .A(n85), .B(n1196), .C(n1195), .D(n1666), .Z(n918) );
  COND2X1 U741 ( .A(n85), .B(n1197), .C(n1196), .D(n1666), .Z(n919) );
  CND2IX1 U758 ( .B(n1687), .A(n1682), .Z(n1199) );
  COND2X1 U798 ( .A(n69), .B(n1222), .C(n1221), .D(n66), .Z(n942) );
  COND2X1 U799 ( .A(n69), .B(n1223), .C(n1222), .D(n66), .Z(n943) );
  COND2X1 U800 ( .A(n69), .B(n1224), .C(n1223), .D(n66), .Z(n944) );
  COND2X1 U801 ( .A(n69), .B(n1225), .C(n1224), .D(n66), .Z(n945) );
  COND2X1 U803 ( .A(n69), .B(n1227), .C(n1226), .D(n66), .Z(n947) );
  COND2X1 U806 ( .A(n69), .B(n1230), .C(n1229), .D(n66), .Z(n950) );
  COND2X1 U809 ( .A(n69), .B(n1233), .C(n1232), .D(n66), .Z(n953) );
  COND2X1 U836 ( .A(n61), .B(n1241), .C(n1240), .D(n58), .Z(n960) );
  COND2X1 U837 ( .A(n61), .B(n1242), .C(n1241), .D(n58), .Z(n961) );
  COND2X1 U838 ( .A(n61), .B(n1243), .C(n1242), .D(n58), .Z(n962) );
  COND2X1 U839 ( .A(n61), .B(n1244), .C(n1243), .D(n58), .Z(n963) );
  COND2X1 U841 ( .A(n61), .B(n1246), .C(n1245), .D(n58), .Z(n965) );
  COND2X1 U842 ( .A(n61), .B(n1247), .C(n1246), .D(n58), .Z(n966) );
  COND2X1 U844 ( .A(n61), .B(n1249), .C(n1248), .D(n58), .Z(n968) );
  COND2X1 U845 ( .A(n61), .B(n1250), .C(n1249), .D(n58), .Z(n969) );
  COND2X1 U847 ( .A(n61), .B(n1252), .C(n1251), .D(n58), .Z(n971) );
  COND2X1 U848 ( .A(n61), .B(n1253), .C(n1252), .D(n58), .Z(n972) );
  COND2X1 U878 ( .A(n53), .B(n1262), .C(n1261), .D(n50), .Z(n980) );
  COND2X1 U879 ( .A(n53), .B(n1263), .C(n1262), .D(n50), .Z(n981) );
  COND2X1 U880 ( .A(n53), .B(n1264), .C(n1263), .D(n50), .Z(n982) );
  COND2X1 U881 ( .A(n53), .B(n1265), .C(n1264), .D(n50), .Z(n983) );
  COND2X1 U883 ( .A(n53), .B(n1267), .C(n1266), .D(n50), .Z(n985) );
  COND2X1 U884 ( .A(n53), .B(n1268), .C(n1267), .D(n50), .Z(n986) );
  COND2X1 U889 ( .A(n53), .B(n1273), .C(n1272), .D(n50), .Z(n991) );
  COND2X1 U890 ( .A(n53), .B(n1274), .C(n1273), .D(n50), .Z(n992) );
  COND2X1 U891 ( .A(n53), .B(n1275), .C(n1274), .D(n50), .Z(n993) );
  COND2X1 U924 ( .A(n44), .B(n1285), .C(n1284), .D(n42), .Z(n1002) );
  COND2X1 U925 ( .A(n44), .B(n1286), .C(n1285), .D(n42), .Z(n1003) );
  COND2X1 U926 ( .A(n44), .B(n1287), .C(n1286), .D(n42), .Z(n1004) );
  COND2X1 U929 ( .A(n44), .B(n1290), .C(n1289), .D(n42), .Z(n1007) );
  COND2X1 U930 ( .A(n44), .B(n1291), .C(n1290), .D(n42), .Z(n1008) );
  COND2X1 U931 ( .A(n44), .B(n1292), .C(n1291), .D(n42), .Z(n1009) );
  COND2X1 U932 ( .A(n44), .B(n1293), .C(n1292), .D(n42), .Z(n1010) );
  COND2X1 U934 ( .A(n44), .B(n1295), .C(n1294), .D(n42), .Z(n1012) );
  COND2X1 U935 ( .A(n44), .B(n1296), .C(n1295), .D(n42), .Z(n1013) );
  COND2X1 U937 ( .A(n44), .B(n1298), .C(n1297), .D(n42), .Z(n1015) );
  COND2X1 U938 ( .A(n44), .B(n1299), .C(n1298), .D(n42), .Z(n1016) );
  COND2X1 U939 ( .A(n44), .B(n1300), .C(n1299), .D(n42), .Z(n1017) );
  COND2X1 U941 ( .A(n44), .B(n1302), .C(n1301), .D(n42), .Z(n1019) );
  CND2IX1 U968 ( .B(n1687), .A(n1709), .Z(n1304) );
  COND2X1 U974 ( .A(n1669), .B(n1310), .C(n1309), .D(n33), .Z(n1026) );
  COND2X1 U975 ( .A(n1669), .B(n1311), .C(n1310), .D(n33), .Z(n1027) );
  COND2X1 U976 ( .A(n36), .B(n1312), .C(n1311), .D(n33), .Z(n1028) );
  COND2X1 U977 ( .A(n36), .B(n1313), .C(n1312), .D(n33), .Z(n1029) );
  COND2X1 U978 ( .A(n1669), .B(n1314), .C(n1313), .D(n33), .Z(n1030) );
  COND2X1 U979 ( .A(n36), .B(n1315), .C(n1314), .D(n33), .Z(n1031) );
  COND2X1 U981 ( .A(n1668), .B(n1317), .C(n1316), .D(n33), .Z(n1033) );
  COND2X1 U982 ( .A(n1669), .B(n1318), .C(n1317), .D(n33), .Z(n1034) );
  COND2X1 U983 ( .A(n1668), .B(n1319), .C(n1318), .D(n33), .Z(n1035) );
  COND2X1 U985 ( .A(n1668), .B(n1321), .C(n1320), .D(n33), .Z(n1037) );
  COND2X1 U988 ( .A(n1669), .B(n1324), .C(n1323), .D(n33), .Z(n1040) );
  COND2X1 U989 ( .A(n1669), .B(n1325), .C(n1324), .D(n33), .Z(n1041) );
  COND2X1 U991 ( .A(n1668), .B(n1327), .C(n1326), .D(n33), .Z(n1043) );
  COND2X1 U1028 ( .A(n27), .B(n1337), .C(n1336), .D(n24), .Z(n1052) );
  COND2X1 U1029 ( .A(n27), .B(n1338), .C(n1337), .D(n24), .Z(n1053) );
  COND2X1 U1030 ( .A(n27), .B(n1339), .C(n1338), .D(n24), .Z(n1054) );
  COND2X1 U1034 ( .A(n27), .B(n1343), .C(n1342), .D(n24), .Z(n1058) );
  COND2X1 U1035 ( .A(n27), .B(n1344), .C(n1343), .D(n24), .Z(n1059) );
  COND2X1 U1037 ( .A(n27), .B(n1346), .C(n1345), .D(n24), .Z(n1061) );
  COND2X1 U1038 ( .A(n27), .B(n1347), .C(n1346), .D(n24), .Z(n1062) );
  COND2X1 U1040 ( .A(n27), .B(n1349), .C(n1348), .D(n24), .Z(n1064) );
  COND2X1 U1042 ( .A(n27), .B(n1351), .C(n1350), .D(n24), .Z(n1066) );
  COND2X1 U1043 ( .A(n27), .B(n1352), .C(n1351), .D(n24), .Z(n1067) );
  COND2X1 U1046 ( .A(n27), .B(n1355), .C(n1354), .D(n24), .Z(n1070) );
  CND2IX1 U1080 ( .B(n1687), .A(n1698), .Z(n1360) );
  COND2X1 U1082 ( .A(n18), .B(n1362), .C(n1661), .D(n1361), .Z(n1076) );
  COND2X1 U1083 ( .A(n18), .B(n1363), .C(n1661), .D(n1362), .Z(n1077) );
  COND2X1 U1084 ( .A(n18), .B(n1364), .C(n1661), .D(n1363), .Z(n1078) );
  COND2X1 U1085 ( .A(n18), .B(n1365), .C(n1661), .D(n1364), .Z(n1079) );
  COND2X1 U1086 ( .A(n18), .B(n1366), .C(n1661), .D(n1365), .Z(n1080) );
  COND2X1 U1087 ( .A(n18), .B(n1367), .C(n1662), .D(n1366), .Z(n1081) );
  COND2X1 U1088 ( .A(n18), .B(n1368), .C(n1661), .D(n1367), .Z(n1082) );
  COND2X1 U1089 ( .A(n18), .B(n1369), .C(n1662), .D(n1368), .Z(n1083) );
  COND2X1 U1090 ( .A(n18), .B(n1370), .C(n1661), .D(n1369), .Z(n1084) );
  COND2X1 U1091 ( .A(n18), .B(n1371), .C(n1661), .D(n1370), .Z(n1085) );
  COND2X1 U1092 ( .A(n18), .B(n1372), .C(n1661), .D(n1371), .Z(n1086) );
  COND2X1 U1093 ( .A(n18), .B(n1373), .C(n1661), .D(n1372), .Z(n1087) );
  COND2X1 U1094 ( .A(n18), .B(n1374), .C(n1662), .D(n1373), .Z(n1088) );
  COND2X1 U1095 ( .A(n18), .B(n1375), .C(n1662), .D(n1374), .Z(n1089) );
  COND2X1 U1096 ( .A(n18), .B(n1376), .C(n1662), .D(n1375), .Z(n1090) );
  COND2X1 U1097 ( .A(n18), .B(n1377), .C(n1662), .D(n1376), .Z(n1091) );
  COND2X1 U1098 ( .A(n18), .B(n1378), .C(n1661), .D(n1377), .Z(n1092) );
  COND2X1 U1099 ( .A(n18), .B(n1379), .C(n1661), .D(n1378), .Z(n1093) );
  COND2X1 U1100 ( .A(n18), .B(n1380), .C(n1662), .D(n1379), .Z(n1094) );
  COND2X1 U1101 ( .A(n18), .B(n1381), .C(n1662), .D(n1380), .Z(n1095) );
  COND2X1 U1102 ( .A(n18), .B(n1382), .C(n1662), .D(n1381), .Z(n1096) );
  COND2X1 U1103 ( .A(n18), .B(n1383), .C(n1662), .D(n1382), .Z(n1097) );
  COND2X1 U1104 ( .A(n18), .B(n1384), .C(n1662), .D(n1383), .Z(n1098) );
  COND2X1 U1105 ( .A(n18), .B(n1385), .C(n1661), .D(n1384), .Z(n1099) );
  COND2X1 U1106 ( .A(n18), .B(n1386), .C(n1662), .D(n1385), .Z(n1100) );
  COND2X1 U1107 ( .A(n18), .B(n1387), .C(n1661), .D(n1386), .Z(n1101) );
  COND2X1 U1108 ( .A(n18), .B(n1388), .C(n1662), .D(n1387), .Z(n1102) );
  COND2X1 U1109 ( .A(n18), .B(n1389), .C(n1661), .D(n1388), .Z(n1103) );
  COND2X1 U1110 ( .A(n1390), .B(n18), .C(n1662), .D(n1389), .Z(n1104) );
  COND2X1 U1144 ( .A(n9), .B(n1393), .C(n6), .D(n1392), .Z(n1106) );
  COND2X1 U1145 ( .A(n9), .B(n1394), .C(n6), .D(n1393), .Z(n1107) );
  COND2X1 U1146 ( .A(n9), .B(n1395), .C(n6), .D(n1394), .Z(n1108) );
  COND2X1 U1147 ( .A(n9), .B(n1396), .C(n6), .D(n1395), .Z(n1109) );
  COND2X1 U1148 ( .A(n9), .B(n1397), .C(n6), .D(n1396), .Z(n1110) );
  COND2X1 U1149 ( .A(n9), .B(n1398), .C(n6), .D(n1397), .Z(n1111) );
  COND2X1 U1150 ( .A(n9), .B(n1399), .C(n6), .D(n1398), .Z(n1112) );
  COND2X1 U1153 ( .A(n9), .B(n1402), .C(n6), .D(n1401), .Z(n1115) );
  COND2X1 U1154 ( .A(n9), .B(n1403), .C(n6), .D(n1402), .Z(n1116) );
  COND2X1 U1155 ( .A(n9), .B(n1404), .C(n6), .D(n1403), .Z(n1117) );
  COND2X1 U1156 ( .A(n9), .B(n1405), .C(n6), .D(n1404), .Z(n1118) );
  COND2X1 U1157 ( .A(n9), .B(n1406), .C(n6), .D(n1405), .Z(n1119) );
  COND2X1 U1158 ( .A(n9), .B(n1407), .C(n6), .D(n1406), .Z(n1120) );
  COND2X1 U1159 ( .A(n9), .B(n1408), .C(n6), .D(n1407), .Z(n1121) );
  COND2X1 U1160 ( .A(n9), .B(n1409), .C(n6), .D(n1408), .Z(n1122) );
  COND2X1 U1161 ( .A(n9), .B(n1410), .C(n6), .D(n1409), .Z(n1123) );
  COND2X1 U1162 ( .A(n9), .B(n1411), .C(n6), .D(n1410), .Z(n1124) );
  COND2X1 U1163 ( .A(n9), .B(n1412), .C(n6), .D(n1411), .Z(n1125) );
  COND2X1 U1164 ( .A(n9), .B(n1413), .C(n6), .D(n1412), .Z(n1126) );
  COND2X1 U1165 ( .A(n9), .B(n1414), .C(n6), .D(n1413), .Z(n1127) );
  COND2X1 U1166 ( .A(n9), .B(n1415), .C(n6), .D(n1414), .Z(n1128) );
  COND2X1 U1167 ( .A(n9), .B(n1416), .C(n6), .D(n1415), .Z(n1129) );
  COND2X1 U1168 ( .A(n9), .B(n1417), .C(n6), .D(n1416), .Z(n1130) );
  COND2X1 U1169 ( .A(n9), .B(n1418), .C(n6), .D(n1417), .Z(n1131) );
  COND2X1 U1170 ( .A(n9), .B(n1419), .C(n6), .D(n1418), .Z(n1132) );
  COND2X1 U1171 ( .A(n9), .B(n1420), .C(n6), .D(n1419), .Z(n1133) );
  COND2X1 U1172 ( .A(n9), .B(n1421), .C(n6), .D(n1420), .Z(n1134) );
  COND2X1 U1173 ( .A(n9), .B(n1422), .C(n6), .D(n1421), .Z(n1135) );
  COND2X1 U1174 ( .A(n1423), .B(n9), .C(n6), .D(n1422), .Z(n1136) );
  CEOX2 U1274 ( .A(a[2]), .B(n1696), .Z(n1457) );
  COND2X1 U1281 ( .A(n1171), .B(n95), .C(n1590), .D(n97), .Z(n854) );
  CIVX1 U1282 ( .A(n891), .Z(n1616) );
  CND2X2 U1283 ( .A(n1445), .B(n105), .Z(n107) );
  CNIVX8 U1284 ( .A(n71), .Z(n1681) );
  CENX1 U1285 ( .A(n1681), .B(n134), .Z(n1207) );
  CENX1 U1286 ( .A(n1681), .B(n136), .Z(n1206) );
  CENX1 U1287 ( .A(n1681), .B(n132), .Z(n1208) );
  CENX1 U1288 ( .A(n1681), .B(n130), .Z(n1209) );
  CENX1 U1289 ( .A(n1681), .B(n146), .Z(n1201) );
  CENXL U1290 ( .A(n1710), .B(n1689), .Z(n1302) );
  CENXL U1291 ( .A(n1710), .B(n152), .Z(n1285) );
  CENXL U1292 ( .A(n1710), .B(n1677), .Z(n1301) );
  CIVXL U1293 ( .A(n223), .Z(n388) );
  CENXL U1294 ( .A(n1686), .B(n1684), .Z(n1170) );
  CENXL U1295 ( .A(n1686), .B(n1683), .Z(n1183) );
  CENXL U1296 ( .A(n1686), .B(n1685), .Z(n1159) );
  CHA1XL U1297 ( .A(n882), .B(n890), .CO(n536), .S(n537) );
  CENX1 U1298 ( .A(n1722), .B(n134), .Z(n1226) );
  CENXL U1299 ( .A(n1695), .B(n138), .Z(n1380) );
  CENXL U1300 ( .A(n1562), .B(n138), .Z(n1413) );
  CENXL U1301 ( .A(n1706), .B(n138), .Z(n1320) );
  CENXL U1302 ( .A(n1718), .B(n138), .Z(n1245) );
  CENXL U1303 ( .A(n1681), .B(n138), .Z(n1205) );
  CND2IX4 U1304 ( .B(n1637), .A(n42), .Z(n44) );
  CENXL U1305 ( .A(n1690), .B(b[30]), .Z(n1393) );
  CENXL U1306 ( .A(n1690), .B(b[29]), .Z(n1394) );
  CENXL U1307 ( .A(n1690), .B(b[28]), .Z(n1395) );
  CENXL U1308 ( .A(n1690), .B(n155), .Z(n1402) );
  CANR1X1 U1309 ( .A(n373), .B(n1655), .C(n370), .Z(n368) );
  CENXL U1310 ( .A(n136), .B(n1684), .Z(n1161) );
  CENXL U1311 ( .A(n1562), .B(n136), .Z(n1414) );
  CENXL U1312 ( .A(n1695), .B(n136), .Z(n1381) );
  CENXL U1313 ( .A(n1706), .B(n136), .Z(n1321) );
  CENXL U1314 ( .A(n1700), .B(n136), .Z(n1350) );
  CENXL U1315 ( .A(n1683), .B(n136), .Z(n1174) );
  CENXL U1316 ( .A(n1716), .B(n136), .Z(n1269) );
  CENXL U1317 ( .A(n1718), .B(n136), .Z(n1246) );
  CENXL U1318 ( .A(n1722), .B(n136), .Z(n1225) );
  CNIVX1 U1319 ( .A(n1018), .Z(n1557) );
  CIVX2 U1320 ( .A(n1564), .Z(n1558) );
  CIVX2 U1321 ( .A(n1558), .Z(n1559) );
  CIVX1 U1322 ( .A(n1558), .Z(n1560) );
  CNIVX1 U1323 ( .A(n1000), .Z(n1561) );
  CENXL U1324 ( .A(n1719), .B(n153), .Z(n1236) );
  CENXL U1325 ( .A(n1690), .B(n153), .Z(n1404) );
  CENXL U1326 ( .A(n1673), .B(n153), .Z(n1259) );
  CENXL U1327 ( .A(n1692), .B(n153), .Z(n1371) );
  CENXL U1328 ( .A(n1698), .B(n153), .Z(n1340) );
  CENXL U1329 ( .A(n132), .B(n1685), .Z(n1152) );
  CENXL U1330 ( .A(n1693), .B(n132), .Z(n1383) );
  CENXL U1331 ( .A(n1690), .B(n132), .Z(n1416) );
  CENXL U1332 ( .A(n1699), .B(n132), .Z(n1352) );
  CENXL U1333 ( .A(n132), .B(n1684), .Z(n1163) );
  CENXL U1334 ( .A(n1704), .B(n132), .Z(n1323) );
  CENXL U1335 ( .A(n1709), .B(n132), .Z(n1296) );
  CENXL U1336 ( .A(n1683), .B(n132), .Z(n1176) );
  CENXL U1337 ( .A(n1718), .B(n132), .Z(n1248) );
  CENXL U1338 ( .A(n1722), .B(n132), .Z(n1227) );
  CENXL U1339 ( .A(n1693), .B(n130), .Z(n1384) );
  CENXL U1340 ( .A(n1699), .B(n130), .Z(n1353) );
  CENXL U1341 ( .A(n130), .B(n1684), .Z(n1164) );
  CENXL U1342 ( .A(n1709), .B(n130), .Z(n1297) );
  CENXL U1343 ( .A(n1704), .B(n130), .Z(n1324) );
  CENXL U1344 ( .A(n1562), .B(n130), .Z(n1417) );
  CENXL U1345 ( .A(n130), .B(n1685), .Z(n1153) );
  CENXL U1346 ( .A(n1715), .B(n130), .Z(n1272) );
  CENXL U1347 ( .A(n1718), .B(n130), .Z(n1249) );
  CENXL U1348 ( .A(n1683), .B(n130), .Z(n1177) );
  CENXL U1349 ( .A(n1704), .B(n134), .Z(n1322) );
  CENXL U1350 ( .A(n1562), .B(n134), .Z(n1415) );
  CENXL U1351 ( .A(n1695), .B(n134), .Z(n1382) );
  CENXL U1352 ( .A(n1683), .B(n134), .Z(n1175) );
  CENXL U1353 ( .A(n1700), .B(n134), .Z(n1351) );
  CENXL U1354 ( .A(n134), .B(n1684), .Z(n1162) );
  CENXL U1355 ( .A(n1709), .B(n134), .Z(n1295) );
  CENXL U1356 ( .A(n1718), .B(n134), .Z(n1247) );
  CENXL U1357 ( .A(n1682), .B(n134), .Z(n1190) );
  CENXL U1358 ( .A(n1683), .B(n140), .Z(n1172) );
  CENXL U1359 ( .A(n1694), .B(n140), .Z(n1379) );
  CENXL U1360 ( .A(n1562), .B(n140), .Z(n1412) );
  CENXL U1361 ( .A(n1706), .B(n140), .Z(n1319) );
  CENXL U1362 ( .A(n1699), .B(n140), .Z(n1348) );
  CENXL U1363 ( .A(n1681), .B(n140), .Z(n1204) );
  CENXL U1364 ( .A(n1718), .B(n140), .Z(n1244) );
  CENXL U1365 ( .A(n1716), .B(n140), .Z(n1267) );
  CENXL U1366 ( .A(n1682), .B(n140), .Z(n1187) );
  CENXL U1367 ( .A(n1722), .B(n140), .Z(n1223) );
  CENXL U1368 ( .A(n1710), .B(n140), .Z(n1292) );
  CENX1 U1369 ( .A(n1719), .B(n152), .Z(n1237) );
  CIVX2 U1370 ( .A(n1618), .Z(n1619) );
  CND2X2 U1371 ( .A(n1450), .B(n74), .Z(n77) );
  CND2X2 U1372 ( .A(n89), .B(n1448), .Z(n91) );
  COND2X1 U1373 ( .A(n1151), .B(n105), .C(n1470), .D(n107), .Z(n852) );
  CNIVX2 U1374 ( .A(n120), .Z(n1688) );
  CNIVX1 U1375 ( .A(n116), .Z(n1686) );
  CND2X1 U1376 ( .A(n1648), .B(n1647), .Z(n245) );
  CENX1 U1377 ( .A(n1698), .B(n146), .Z(n1345) );
  CENX1 U1378 ( .A(n1681), .B(n1677), .Z(n1213) );
  CENX1 U1379 ( .A(n1681), .B(n1678), .Z(n1212) );
  CNR2X1 U1380 ( .A(n69), .B(n1228), .Z(n1605) );
  CENX1 U1381 ( .A(n1677), .B(n1682), .Z(n1196) );
  CENX1 U1382 ( .A(n1681), .B(n1679), .Z(n1211) );
  CENX1 U1383 ( .A(n1721), .B(n130), .Z(n1228) );
  CENX1 U1384 ( .A(n1701), .B(n148), .Z(n1344) );
  CENX1 U1385 ( .A(n1678), .B(n1683), .Z(n1180) );
  CENX1 U1386 ( .A(n1682), .B(n130), .Z(n1192) );
  CENX1 U1387 ( .A(n1687), .B(n1719), .Z(n1255) );
  CENX1 U1388 ( .A(n1718), .B(n1688), .Z(n1254) );
  CENX1 U1389 ( .A(n1687), .B(n1722), .Z(n1234) );
  CENX1 U1390 ( .A(n1560), .B(n148), .Z(n1408) );
  CENX1 U1391 ( .A(n1560), .B(n146), .Z(n1409) );
  CENX1 U1392 ( .A(n1718), .B(n1678), .Z(n1252) );
  CENX1 U1393 ( .A(n1718), .B(n1677), .Z(n1253) );
  CENX1 U1394 ( .A(n1700), .B(n138), .Z(n1349) );
  CENX1 U1395 ( .A(n1560), .B(n150), .Z(n1407) );
  CENX1 U1396 ( .A(n1718), .B(n1680), .Z(n1250) );
  CENX1 U1397 ( .A(n1718), .B(n1679), .Z(n1251) );
  CENX1 U1398 ( .A(n1688), .B(n1681), .Z(n1214) );
  CENX1 U1399 ( .A(n1687), .B(n1681), .Z(n1215) );
  CENX1 U1400 ( .A(n1673), .B(n132), .Z(n1271) );
  CENX1 U1401 ( .A(n1560), .B(n151), .Z(n1406) );
  CENX1 U1402 ( .A(n1711), .B(n138), .Z(n1293) );
  CENX1 U1403 ( .A(n1716), .B(n138), .Z(n1268) );
  CENX1 U1404 ( .A(n1690), .B(n156), .Z(n1401) );
  CENX1 U1405 ( .A(n1681), .B(n1680), .Z(n1210) );
  CENX1 U1406 ( .A(n1688), .B(n1683), .Z(n1182) );
  CENX1 U1407 ( .A(n1677), .B(n1683), .Z(n1181) );
  CENX1 U1408 ( .A(n1690), .B(n154), .Z(n1403) );
  CIVX2 U1409 ( .A(n48), .Z(n1717) );
  CENX1 U1410 ( .A(n1721), .B(n142), .Z(n1222) );
  CENX1 U1411 ( .A(n1719), .B(n146), .Z(n1241) );
  COND2X1 U1412 ( .A(n1160), .B(n1609), .C(n1471), .D(n102), .Z(n853) );
  CENX1 U1413 ( .A(n1673), .B(n146), .Z(n1264) );
  CENX1 U1414 ( .A(n1716), .B(n148), .Z(n1263) );
  CENX1 U1415 ( .A(n1680), .B(n1683), .Z(n1178) );
  CENX1 U1416 ( .A(n1679), .B(n1683), .Z(n1179) );
  CENX1 U1417 ( .A(n1718), .B(n142), .Z(n1243) );
  CENX1 U1418 ( .A(n1719), .B(n148), .Z(n1240) );
  CENX1 U1419 ( .A(n1719), .B(n150), .Z(n1239) );
  CENX1 U1420 ( .A(n1681), .B(n142), .Z(n1203) );
  CENX1 U1421 ( .A(n1690), .B(b[26]), .Z(n1397) );
  CENX1 U1422 ( .A(n1716), .B(n150), .Z(n1262) );
  CENX1 U1423 ( .A(n1560), .B(n142), .Z(n1411) );
  CENX1 U1424 ( .A(n1686), .B(n1702), .Z(n1359) );
  CNIVX3 U1425 ( .A(n122), .Z(n1677) );
  CNIVX2 U1426 ( .A(n126), .Z(n1679) );
  CNIVX2 U1427 ( .A(n128), .Z(n1680) );
  CENX1 U1428 ( .A(n1688), .B(n109), .Z(n1142) );
  CENX1 U1429 ( .A(n1719), .B(n151), .Z(n1238) );
  CIVX2 U1430 ( .A(n1659), .Z(n42) );
  CNIVX2 U1431 ( .A(n124), .Z(n1678) );
  CENX1 U1432 ( .A(n1677), .B(n109), .Z(n1141) );
  CND2X1 U1433 ( .A(n1601), .B(n1602), .Z(n1449) );
  CND2X1 U1434 ( .A(n1599), .B(n1682), .Z(n1602) );
  CND3X1 U1435 ( .A(n1574), .B(n1575), .C(n1576), .Z(n528) );
  CENX1 U1436 ( .A(n1694), .B(n1688), .Z(n1389) );
  CENX1 U1437 ( .A(n1694), .B(b[29]), .Z(n1361) );
  CNIVX1 U1438 ( .A(n15), .Z(n1660) );
  CENX1 U1439 ( .A(n1681), .B(n148), .Z(n1200) );
  CENX1 U1440 ( .A(n1722), .B(n151), .Z(n1217) );
  CANR1X1 U1441 ( .A(n257), .B(n1648), .C(n248), .Z(n246) );
  CNR2X1 U1442 ( .A(n1570), .B(n512), .Z(n218) );
  CNIVX2 U1443 ( .A(n116), .Z(n1687) );
  COND1XL U1444 ( .A(n376), .B(n374), .C(n375), .Z(n373) );
  CENX1 U1445 ( .A(n1686), .B(n1560), .Z(n1423) );
  CANR1X1 U1446 ( .A(n275), .B(n1643), .C(n268), .Z(n262) );
  CNR2X1 U1447 ( .A(n513), .B(n538), .Z(n223) );
  CENX1 U1448 ( .A(n271), .B(n175), .Z(product[22]) );
  CIVX2 U1449 ( .A(n242), .Z(n241) );
  CFA1XL U1450 ( .A(n1130), .B(n1100), .CI(n1072), .CO(n834), .S(n835) );
  CIVX1 U1451 ( .A(n216), .Z(n1597) );
  CENX1 U1452 ( .A(n1710), .B(n1678), .Z(n1300) );
  CIVX3 U1453 ( .A(n1713), .Z(n1710) );
  CFA1XL U1454 ( .A(n959), .B(n1079), .CI(n1051), .CO(n504), .S(n505) );
  CIVX4 U1455 ( .A(n1636), .Z(n24) );
  CEOX2 U1456 ( .A(n1694), .B(a[4]), .Z(n1636) );
  CENXL U1457 ( .A(n1686), .B(n1696), .Z(n1390) );
  CNR2IX1 U1458 ( .B(n1687), .A(n110), .Z(n871) );
  CIVX2 U1459 ( .A(n30), .Z(n1708) );
  CIVX2 U1460 ( .A(n1708), .Z(n1704) );
  CNIVX2 U1461 ( .A(n1691), .Z(n1562) );
  CIVDX1 U1462 ( .A(n3), .Z0(n1563), .Z1(n1564) );
  CIVX2 U1463 ( .A(n12), .Z(n1697) );
  CIVX1 U1464 ( .A(n1697), .Z(n1693) );
  COND2X1 U1465 ( .A(n85), .B(n1187), .C(n1186), .D(n1666), .Z(n909) );
  CIVX2 U1466 ( .A(n74), .Z(n1618) );
  CIVX2 U1467 ( .A(n1684), .Z(n1590) );
  COAN1X1 U1468 ( .A(n330), .B(n313), .C(n314), .Z(n1565) );
  COR2X1 U1469 ( .A(n1136), .B(n865), .Z(n1566) );
  CANR1X1 U1470 ( .A(n1640), .B(n213), .C(n210), .Z(n208) );
  COND2XL U1471 ( .A(n53), .B(n1276), .C(n1275), .D(n50), .Z(n994) );
  CIVXL U1472 ( .A(n234), .Z(n389) );
  CENX1 U1473 ( .A(n1686), .B(n1673), .Z(n1278) );
  CENX1 U1474 ( .A(n1716), .B(n151), .Z(n1261) );
  COND2XL U1475 ( .A(n1234), .B(n69), .C(n1233), .D(n66), .Z(n954) );
  CENXL U1476 ( .A(n241), .B(n172), .Z(product[25]) );
  CENXL U1477 ( .A(n1567), .B(n227), .Z(product[27]) );
  CAN2X1 U1478 ( .A(n388), .B(n226), .Z(n1567) );
  CND2X1 U1479 ( .A(a[22]), .B(n1590), .Z(n1591) );
  CENXL U1480 ( .A(n1568), .B(n236), .Z(product[26]) );
  CAN2XL U1481 ( .A(n389), .B(n235), .Z(n1568) );
  CND2X1 U1482 ( .A(n1624), .B(n1625), .Z(n1627) );
  CIVX2 U1483 ( .A(n1718), .Z(n1624) );
  CND2X4 U1484 ( .A(n95), .B(n1447), .Z(n97) );
  COND2XL U1485 ( .A(n44), .B(n1281), .C(n1280), .D(n42), .Z(n998) );
  COND2XL U1486 ( .A(n44), .B(n1282), .C(n1281), .D(n42), .Z(n999) );
  COND2XL U1487 ( .A(n44), .B(n1294), .C(n1293), .D(n42), .Z(n1011) );
  COND2XL U1488 ( .A(n44), .B(n1713), .C(n42), .D(n1304), .Z(n861) );
  COND2XL U1489 ( .A(n1303), .B(n44), .C(n1302), .D(n42), .Z(n1020) );
  COND2XL U1490 ( .A(n44), .B(n1284), .C(n1283), .D(n42), .Z(n1001) );
  COND2XL U1491 ( .A(n44), .B(n1283), .C(n1282), .D(n42), .Z(n1000) );
  COND2XL U1492 ( .A(n44), .B(n1301), .C(n1300), .D(n42), .Z(n1018) );
  COND2XL U1493 ( .A(n44), .B(n1288), .C(n1287), .D(n42), .Z(n1005) );
  COND2XL U1494 ( .A(n44), .B(n1297), .C(n1296), .D(n42), .Z(n1014) );
  CENXL U1495 ( .A(n1569), .B(n199), .Z(product[31]) );
  CAN2X1 U1496 ( .A(n1653), .B(n198), .Z(n1569) );
  CND2X1 U1497 ( .A(n1455), .B(n33), .Z(n36) );
  CND2X1 U1498 ( .A(n1455), .B(n33), .Z(n1668) );
  CEOX2 U1499 ( .A(a[6]), .B(n1704), .Z(n1455) );
  COND2X1 U1500 ( .A(n44), .B(n1289), .C(n1288), .D(n42), .Z(n1006) );
  CENX1 U1501 ( .A(n1673), .B(n142), .Z(n1266) );
  CFA1XL U1502 ( .A(n949), .B(n1087), .CI(n1009), .CO(n684), .S(n685) );
  CHA1XL U1503 ( .A(n860), .B(n996), .CO(n808), .S(n809) );
  CIVX1 U1504 ( .A(n330), .Z(n329) );
  COND2X1 U1505 ( .A(n61), .B(n1248), .C(n1247), .D(n58), .Z(n967) );
  CFA1XL U1506 ( .A(n1021), .B(n1129), .CI(n1045), .CO(n830), .S(n831) );
  COND1X1 U1507 ( .A(n299), .B(n295), .C(n296), .Z(n294) );
  COND2XL U1508 ( .A(n69), .B(n1232), .C(n1231), .D(n66), .Z(n952) );
  COND2XL U1509 ( .A(n69), .B(n1220), .C(n1219), .D(n66), .Z(n940) );
  COND2XL U1510 ( .A(n69), .B(n1229), .C(n1228), .D(n66), .Z(n949) );
  COND2XL U1511 ( .A(n69), .B(n1221), .C(n1220), .D(n66), .Z(n941) );
  CNR2IXL U1512 ( .B(n1687), .A(n66), .Z(n955) );
  CEO3X1 U1513 ( .A(n491), .B(n489), .C(n514), .Z(n1570) );
  CEO3XL U1514 ( .A(n491), .B(n489), .C(n514), .Z(n1571) );
  CFA1XL U1515 ( .A(n491), .B(n489), .CI(n514), .CO(n486), .S(n487) );
  CENX2 U1516 ( .A(n1681), .B(a[18]), .Z(n1666) );
  CENX1 U1517 ( .A(n1690), .B(b[24]), .Z(n1399) );
  CENX1 U1518 ( .A(n1690), .B(b[25]), .Z(n1398) );
  CIVX2 U1519 ( .A(n229), .Z(n1596) );
  CNR2XL U1520 ( .A(n234), .B(n239), .Z(n228) );
  COND2X1 U1521 ( .A(n1668), .B(n1309), .C(n1308), .D(n33), .Z(n1025) );
  CND2IXL U1522 ( .B(n1687), .A(n1683), .Z(n1184) );
  CENXL U1523 ( .A(n1683), .B(n138), .Z(n1173) );
  CEOX1 U1524 ( .A(a[20]), .B(n1683), .Z(n1448) );
  CND2X1 U1525 ( .A(n1628), .B(n1629), .Z(n1631) );
  COND2X1 U1526 ( .A(n77), .B(n1209), .C(n1208), .D(n1619), .Z(n930) );
  CIVX2 U1527 ( .A(n1717), .Z(n1716) );
  CIVX1 U1528 ( .A(n1717), .Z(n1673) );
  CIVXL U1529 ( .A(n262), .Z(n264) );
  CENXL U1530 ( .A(n1572), .B(n636), .Z(n613) );
  CENXL U1531 ( .A(n638), .B(n619), .Z(n1572) );
  COND2X1 U1532 ( .A(n85), .B(n1191), .C(n1190), .D(n1666), .Z(n913) );
  COND1X1 U1533 ( .A(n262), .B(n245), .C(n246), .Z(n244) );
  CIVXL U1534 ( .A(n279), .Z(n278) );
  CIVX2 U1535 ( .A(n1664), .Z(n1690) );
  CIVX4 U1536 ( .A(n1717), .Z(n1715) );
  COND2X1 U1537 ( .A(n1669), .B(n1323), .C(n1322), .D(n33), .Z(n1039) );
  COND1XL U1538 ( .A(n328), .B(n322), .C(n323), .Z(n321) );
  CIVX1 U1539 ( .A(n322), .Z(n401) );
  CFA1X1 U1540 ( .A(n916), .B(n964), .CI(n1030), .CO(n624), .S(n625) );
  CEOX2 U1541 ( .A(a[14]), .B(n1722), .Z(n1451) );
  CIVX2 U1542 ( .A(n1697), .Z(n1694) );
  COND2X1 U1543 ( .A(n97), .B(n1168), .C(n95), .D(n1167), .Z(n892) );
  COND2X1 U1544 ( .A(n97), .B(n1167), .C(n95), .D(n1166), .Z(n891) );
  COND2XL U1545 ( .A(n1170), .B(n97), .C(n95), .D(n1169), .Z(n894) );
  CEOX2 U1546 ( .A(n30), .B(a[8]), .Z(n1659) );
  CNR2IX1 U1547 ( .B(n1687), .A(n1619), .Z(n937) );
  COND1X1 U1548 ( .A(n280), .B(n292), .C(n281), .Z(n279) );
  CFA1XL U1549 ( .A(n958), .B(n1050), .CI(n1078), .CO(n476), .S(n477) );
  CIVX4 U1550 ( .A(n1720), .Z(n1718) );
  CIVX3 U1551 ( .A(n55), .Z(n1720) );
  CEOX2 U1552 ( .A(a[10]), .B(n1716), .Z(n1453) );
  CEOX1 U1553 ( .A(n602), .B(n583), .Z(n1586) );
  CNR2X1 U1554 ( .A(n223), .B(n218), .Z(n216) );
  CANR1X1 U1555 ( .A(n221), .B(n241), .C(n222), .Z(n220) );
  COND1X1 U1556 ( .A(n226), .B(n218), .C(n219), .Z(n217) );
  CND2XL U1557 ( .A(n513), .B(n538), .Z(n226) );
  CNIVX1 U1558 ( .A(n1056), .Z(n1573) );
  COND2X1 U1559 ( .A(n77), .B(n1208), .C(n1207), .D(n1619), .Z(n929) );
  CND2XL U1560 ( .A(n1648), .B(n250), .Z(n173) );
  CENXL U1561 ( .A(n1690), .B(b[27]), .Z(n1396) );
  CENX1 U1562 ( .A(n1711), .B(n150), .Z(n1287) );
  CIVX1 U1563 ( .A(n1714), .Z(n1711) );
  CIVX2 U1564 ( .A(n39), .Z(n1714) );
  CND2IXL U1565 ( .B(n1687), .A(n1716), .Z(n1279) );
  CENXL U1566 ( .A(n1673), .B(n152), .Z(n1260) );
  CIVX2 U1567 ( .A(n21), .Z(n1703) );
  CND2IXL U1568 ( .B(n1687), .A(n1719), .Z(n1256) );
  CEOX2 U1569 ( .A(a[12]), .B(n1719), .Z(n1452) );
  COND2XL U1570 ( .A(n1668), .B(n1329), .C(n1328), .D(n33), .Z(n1045) );
  COND2XL U1571 ( .A(n1669), .B(n1316), .C(n1315), .D(n33), .Z(n1032) );
  COND2X1 U1572 ( .A(n9), .B(n1401), .C(n6), .D(n1400), .Z(n1114) );
  CANR1X1 U1573 ( .A(n348), .B(n1652), .C(n343), .Z(n341) );
  CNR2X2 U1574 ( .A(n707), .B(n722), .Z(n295) );
  COND2X1 U1575 ( .A(n61), .B(n1251), .C(n1250), .D(n58), .Z(n970) );
  CND2IXL U1576 ( .B(n1687), .A(n1681), .Z(n1216) );
  CND2X2 U1577 ( .A(n1449), .B(n82), .Z(n85) );
  CND2X1 U1578 ( .A(n1718), .B(a[14]), .Z(n1626) );
  COND2X1 U1579 ( .A(n9), .B(n1400), .C(n6), .D(n1399), .Z(n1113) );
  CEO3X2 U1580 ( .A(n1026), .B(n1080), .C(n1052), .Z(n529) );
  CND2X1 U1581 ( .A(n1026), .B(n1052), .Z(n1574) );
  CND2X1 U1582 ( .A(n1080), .B(n1026), .Z(n1575) );
  CND2X1 U1583 ( .A(n1052), .B(n1080), .Z(n1576) );
  CENX4 U1584 ( .A(n1682), .B(a[20]), .Z(n89) );
  CNIVX16 U1585 ( .A(n79), .Z(n1682) );
  CIVX2 U1586 ( .A(n1682), .Z(n1600) );
  COND2XL U1587 ( .A(n61), .B(n1237), .C(n1236), .D(n58), .Z(n956) );
  COND2XL U1588 ( .A(n61), .B(n1238), .C(n1237), .D(n58), .Z(n957) );
  COND2XL U1589 ( .A(n61), .B(n1240), .C(n1239), .D(n58), .Z(n959) );
  COND2XL U1590 ( .A(n61), .B(n1239), .C(n1238), .D(n58), .Z(n958) );
  COND2XL U1591 ( .A(n1255), .B(n61), .C(n1254), .D(n58), .Z(n974) );
  COND2XL U1592 ( .A(n61), .B(n1245), .C(n1244), .D(n58), .Z(n964) );
  COND2X1 U1593 ( .A(n61), .B(n1254), .C(n1253), .D(n58), .Z(n973) );
  CND2X4 U1594 ( .A(n1453), .B(n50), .Z(n53) );
  COND2X1 U1595 ( .A(n53), .B(n1259), .C(n1258), .D(n50), .Z(n977) );
  CENXL U1596 ( .A(n1673), .B(n154), .Z(n1258) );
  CENX1 U1597 ( .A(a[4]), .B(n1702), .Z(n1635) );
  CIVX1 U1598 ( .A(n1703), .Z(n1702) );
  CANR1X1 U1599 ( .A(n288), .B(n1646), .C(n283), .Z(n281) );
  CIVXL U1600 ( .A(n292), .Z(n291) );
  CFA1X1 U1601 ( .A(n1039), .B(n788), .CI(n1065), .CO(n772), .S(n773) );
  COND2X1 U1602 ( .A(n53), .B(n1266), .C(n1265), .D(n50), .Z(n984) );
  COND1X1 U1603 ( .A(n368), .B(n366), .C(n367), .Z(n365) );
  COND1X1 U1604 ( .A(n240), .B(n234), .C(n235), .Z(n229) );
  CND2X2 U1605 ( .A(n563), .B(n586), .Z(n240) );
  CNR2IX1 U1606 ( .B(n1687), .A(n1609), .Z(n885) );
  CNR2XL U1607 ( .A(n27), .B(n1345), .Z(n1577) );
  CNR2XL U1608 ( .A(n1344), .B(n24), .Z(n1578) );
  COR2X1 U1609 ( .A(n1577), .B(n1578), .Z(n1060) );
  CEOX1 U1610 ( .A(n1013), .B(n1121), .Z(n1579) );
  CEOX1 U1611 ( .A(n1579), .B(n1037), .Z(n747) );
  CND2XL U1612 ( .A(n1037), .B(n1121), .Z(n1580) );
  CND2X1 U1613 ( .A(n1037), .B(n1013), .Z(n1581) );
  CND2XL U1614 ( .A(n1121), .B(n1013), .Z(n1582) );
  CND3X1 U1615 ( .A(n1580), .B(n1581), .C(n1582), .Z(n746) );
  CND2XL U1616 ( .A(a[26]), .B(n1470), .Z(n1584) );
  CND2X1 U1617 ( .A(n1583), .B(n104), .Z(n1585) );
  CND2X1 U1618 ( .A(n1584), .B(n1585), .Z(n1445) );
  CIVXL U1619 ( .A(a[26]), .Z(n1583) );
  CEOX2 U1620 ( .A(n1586), .B(n600), .Z(n573) );
  CND2XL U1621 ( .A(n583), .B(n600), .Z(n1587) );
  CND2X1 U1622 ( .A(n600), .B(n602), .Z(n1588) );
  CND2XL U1623 ( .A(n583), .B(n602), .Z(n1589) );
  CND3X1 U1624 ( .A(n1587), .B(n1588), .C(n1589), .Z(n572) );
  CND2XL U1625 ( .A(n1629), .B(n1684), .Z(n1592) );
  CND2X1 U1626 ( .A(n1591), .B(n1592), .Z(n1447) );
  CND2X1 U1627 ( .A(n636), .B(n619), .Z(n1593) );
  CND2X1 U1628 ( .A(n636), .B(n638), .Z(n1594) );
  CND2X1 U1629 ( .A(n619), .B(n638), .Z(n1595) );
  CND3X2 U1630 ( .A(n1593), .B(n1594), .C(n1595), .Z(n612) );
  CND3XL U1631 ( .A(n1674), .B(n1675), .C(n1676), .Z(n638) );
  CNR2X2 U1632 ( .A(n1596), .B(n1597), .Z(n1598) );
  CNR2X2 U1633 ( .A(n1598), .B(n217), .Z(n215) );
  CND2X2 U1634 ( .A(a[18]), .B(n1600), .Z(n1601) );
  CIVX1 U1635 ( .A(a[18]), .Z(n1599) );
  COR2XL U1636 ( .A(n53), .B(n1272), .Z(n1603) );
  COR2XL U1637 ( .A(n1271), .B(n50), .Z(n1604) );
  CND2X1 U1638 ( .A(n1603), .B(n1604), .Z(n990) );
  CNR2XL U1639 ( .A(n1227), .B(n66), .Z(n1606) );
  COR2X1 U1640 ( .A(n1605), .B(n1606), .Z(n948) );
  CND2X4 U1641 ( .A(n1451), .B(n66), .Z(n69) );
  CND2X4 U1642 ( .A(n1626), .B(n1627), .Z(n66) );
  CNIVX4 U1643 ( .A(n87), .Z(n1683) );
  CIVX2 U1644 ( .A(n100), .Z(n1607) );
  CIVX2 U1645 ( .A(n1607), .Z(n1608) );
  CIVX2 U1646 ( .A(n1607), .Z(n1609) );
  CIVXL U1647 ( .A(n917), .Z(n1610) );
  CIVX1 U1648 ( .A(n1610), .Z(n1611) );
  CIVXL U1649 ( .A(n920), .Z(n1612) );
  CIVX1 U1650 ( .A(n1612), .Z(n1613) );
  COND2XL U1651 ( .A(n27), .B(n1333), .C(n1332), .D(n24), .Z(n1048) );
  COND2XL U1652 ( .A(n27), .B(n1334), .C(n1333), .D(n24), .Z(n1049) );
  COND2XL U1653 ( .A(n27), .B(n1356), .C(n1355), .D(n24), .Z(n1071) );
  COND2XL U1654 ( .A(n27), .B(n1354), .C(n1353), .D(n24), .Z(n1069) );
  COND2XL U1655 ( .A(n27), .B(n1353), .C(n1352), .D(n24), .Z(n1068) );
  COND2XL U1656 ( .A(n27), .B(n1357), .C(n1356), .D(n24), .Z(n1072) );
  COND2XL U1657 ( .A(n27), .B(n1341), .C(n1340), .D(n24), .Z(n1056) );
  COND2XL U1658 ( .A(n27), .B(n1336), .C(n1335), .D(n24), .Z(n1051) );
  COND2XL U1659 ( .A(n27), .B(n1335), .C(n1334), .D(n24), .Z(n1050) );
  COND2XL U1660 ( .A(n27), .B(n1350), .C(n1349), .D(n24), .Z(n1065) );
  COND2XL U1661 ( .A(n1359), .B(n27), .C(n1358), .D(n24), .Z(n1074) );
  COND2X1 U1662 ( .A(n27), .B(n1340), .C(n1339), .D(n24), .Z(n1055) );
  COND1X1 U1663 ( .A(n214), .B(n242), .C(n215), .Z(n213) );
  CNR2X1 U1664 ( .A(n245), .B(n261), .Z(n243) );
  CENXL U1665 ( .A(n1682), .B(n144), .Z(n1185) );
  CENXL U1666 ( .A(n1707), .B(n144), .Z(n1317) );
  CENXL U1667 ( .A(n1560), .B(n144), .Z(n1410) );
  CENXL U1668 ( .A(n1696), .B(n144), .Z(n1377) );
  CENXL U1669 ( .A(n1719), .B(n144), .Z(n1242) );
  CENXL U1670 ( .A(n1698), .B(n144), .Z(n1346) );
  CENXL U1671 ( .A(n1723), .B(n144), .Z(n1221) );
  CENXL U1672 ( .A(n1681), .B(n144), .Z(n1202) );
  CENXL U1673 ( .A(n1715), .B(n144), .Z(n1265) );
  CENXL U1674 ( .A(n1710), .B(n144), .Z(n1290) );
  CANR1X1 U1675 ( .A(n1639), .B(n213), .C(n1638), .Z(n199) );
  CIVXL U1676 ( .A(n915), .Z(n1614) );
  CIVX2 U1677 ( .A(n1614), .Z(n1615) );
  CND2X4 U1678 ( .A(n1452), .B(n58), .Z(n61) );
  CIVX1 U1679 ( .A(n1616), .Z(n1617) );
  CEOX2 U1680 ( .A(a[16]), .B(n1681), .Z(n1450) );
  CIVX4 U1681 ( .A(n1658), .Z(n33) );
  CEOX2 U1682 ( .A(n1700), .B(a[6]), .Z(n1658) );
  CENXL U1683 ( .A(n1704), .B(b[25]), .Z(n1305) );
  CENXL U1684 ( .A(n1698), .B(b[25]), .Z(n1334) );
  CENXL U1685 ( .A(n1693), .B(b[25]), .Z(n1365) );
  CIVXL U1686 ( .A(n352), .Z(n351) );
  CENXL U1687 ( .A(n1715), .B(n134), .Z(n1270) );
  CND2X2 U1688 ( .A(n1455), .B(n33), .Z(n1669) );
  COND2XL U1689 ( .A(n85), .B(n1186), .C(n1185), .D(n1666), .Z(n908) );
  COND2XL U1690 ( .A(n85), .B(n1189), .C(n1188), .D(n1666), .Z(n911) );
  COND2XL U1691 ( .A(n85), .B(n1188), .C(n1187), .D(n1666), .Z(n910) );
  COND2XL U1692 ( .A(n85), .B(n1194), .C(n1193), .D(n1666), .Z(n916) );
  COND2XL U1693 ( .A(n85), .B(n1193), .C(n1192), .D(n1666), .Z(n915) );
  COND2XL U1694 ( .A(n1198), .B(n85), .C(n1666), .D(n1197), .Z(n920) );
  COND2XL U1695 ( .A(n85), .B(n1195), .C(n1194), .D(n1666), .Z(n917) );
  CENX2 U1696 ( .A(n1685), .B(a[26]), .Z(n105) );
  CND2IXL U1697 ( .B(n1687), .A(n109), .Z(n1144) );
  CND2XL U1698 ( .A(n1690), .B(n157), .Z(n1622) );
  CND2XL U1699 ( .A(n1620), .B(n1621), .Z(n1623) );
  CND2X1 U1700 ( .A(n1622), .B(n1623), .Z(n1400) );
  CIVXL U1701 ( .A(n1690), .Z(n1620) );
  CIVXL U1702 ( .A(n157), .Z(n1621) );
  CANR1X2 U1703 ( .A(n243), .B(n279), .C(n244), .Z(n242) );
  CIVXL U1704 ( .A(a[14]), .Z(n1625) );
  COND2XL U1705 ( .A(n69), .B(n1218), .C(n1217), .D(n66), .Z(n938) );
  COND2XL U1706 ( .A(n69), .B(n1724), .C(n66), .D(n1235), .Z(n858) );
  COND2XL U1707 ( .A(n69), .B(n1219), .C(n1218), .D(n66), .Z(n939) );
  CIVXL U1708 ( .A(n1685), .Z(n1471) );
  COND2XL U1709 ( .A(n102), .B(n1157), .C(n1609), .D(n1156), .Z(n882) );
  COND2XL U1710 ( .A(n102), .B(n1155), .C(n1609), .D(n1154), .Z(n880) );
  CENXL U1711 ( .A(n1663), .B(n208), .Z(product[30]) );
  CND2XL U1712 ( .A(n1683), .B(a[22]), .Z(n1630) );
  CND2X2 U1713 ( .A(n1630), .B(n1631), .Z(n95) );
  CIVXL U1714 ( .A(n1683), .Z(n1628) );
  CIVXL U1715 ( .A(a[22]), .Z(n1629) );
  COND2XL U1716 ( .A(n97), .B(n1162), .C(n1161), .D(n95), .Z(n886) );
  COND2X1 U1717 ( .A(n97), .B(n1169), .C(n95), .D(n1168), .Z(n893) );
  COND2XL U1718 ( .A(n97), .B(n1166), .C(n95), .D(n1165), .Z(n890) );
  COND2XL U1719 ( .A(n97), .B(n1164), .C(n1163), .D(n95), .Z(n888) );
  COND1X1 U1720 ( .A(n352), .B(n340), .C(n341), .Z(n339) );
  CANR1X1 U1721 ( .A(n1645), .B(n321), .C(n316), .Z(n314) );
  CNR2XL U1722 ( .A(n322), .B(n327), .Z(n320) );
  CND2XL U1723 ( .A(n849), .B(n1104), .Z(n375) );
  CIVX2 U1724 ( .A(n1724), .Z(n1721) );
  CND2X1 U1725 ( .A(n1643), .B(n394), .Z(n261) );
  CNR2X1 U1726 ( .A(n651), .B(n670), .Z(n272) );
  CANR1XL U1727 ( .A(n1650), .B(n357), .C(n354), .Z(n352) );
  CANR1XL U1728 ( .A(n365), .B(n1654), .C(n362), .Z(n360) );
  COR2X1 U1729 ( .A(n819), .B(n826), .Z(n1651) );
  CEO3X1 U1730 ( .A(n452), .B(n450), .C(n448), .Z(n422) );
  CIVX1 U1731 ( .A(n1563), .Z(n1691) );
  CNR2IX1 U1732 ( .B(n1687), .A(n114), .Z(n867) );
  COND2X1 U1733 ( .A(n69), .B(n1231), .C(n1230), .D(n66), .Z(n951) );
  CEO3X1 U1734 ( .A(n428), .B(n427), .C(n426), .Z(n421) );
  CEO3X1 U1735 ( .A(n896), .B(n922), .C(n976), .Z(n427) );
  CENX1 U1736 ( .A(n1684), .B(a[24]), .Z(n100) );
  CENX1 U1737 ( .A(n1673), .B(n155), .Z(n1257) );
  CENX1 U1738 ( .A(n1707), .B(n150), .Z(n1314) );
  CENX1 U1739 ( .A(n1701), .B(n150), .Z(n1343) );
  CENX1 U1740 ( .A(n1723), .B(n150), .Z(n1218) );
  CENX1 U1741 ( .A(n1693), .B(n150), .Z(n1374) );
  CEOXL U1742 ( .A(n1632), .B(n213), .Z(product[29]) );
  CAN2XL U1743 ( .A(n1640), .B(n212), .Z(n1632) );
  CND2XL U1744 ( .A(n390), .B(n240), .Z(n172) );
  CAN2XL U1745 ( .A(n1641), .B(n1640), .Z(n1639) );
  CANR1X1 U1746 ( .A(n312), .B(n293), .C(n294), .Z(n292) );
  CNR2XL U1747 ( .A(n295), .B(n298), .Z(n293) );
  CEOXL U1748 ( .A(n169), .B(n220), .Z(product[28]) );
  CIVX1 U1749 ( .A(n273), .Z(n275) );
  CANR1X1 U1750 ( .A(n308), .B(n1642), .C(n301), .Z(n299) );
  CIVX1 U1751 ( .A(n303), .Z(n301) );
  CND2XL U1752 ( .A(n1645), .B(n318), .Z(n182) );
  CEOXL U1753 ( .A(n182), .B(n319), .Z(product[15]) );
  CEOXL U1754 ( .A(n177), .B(n286), .Z(product[20]) );
  CND2XL U1755 ( .A(n1646), .B(n285), .Z(n177) );
  CEOXL U1756 ( .A(n176), .B(n278), .Z(product[21]) );
  CND2XL U1757 ( .A(n394), .B(n273), .Z(n176) );
  CEOXL U1758 ( .A(n183), .B(n324), .Z(product[14]) );
  CEOXL U1759 ( .A(n181), .B(n1565), .Z(product[16]) );
  CND2XL U1760 ( .A(n399), .B(n306), .Z(n181) );
  CND2XL U1761 ( .A(n1644), .B(n290), .Z(n178) );
  CND2XL U1762 ( .A(n539), .B(n562), .Z(n235) );
  CND2XL U1763 ( .A(n399), .B(n1642), .Z(n298) );
  CND2XL U1764 ( .A(n1571), .B(n512), .Z(n219) );
  CANR1X1 U1765 ( .A(n331), .B(n339), .C(n332), .Z(n330) );
  CNR2XL U1766 ( .A(n333), .B(n336), .Z(n331) );
  CND2XL U1767 ( .A(n767), .B(n778), .Z(n323) );
  CND2XL U1768 ( .A(n1652), .B(n345), .Z(n187) );
  CND2XL U1769 ( .A(n404), .B(n337), .Z(n186) );
  CND2XL U1770 ( .A(n402), .B(n328), .Z(n184) );
  CND2XL U1771 ( .A(n1650), .B(n356), .Z(n189) );
  CND2XL U1772 ( .A(n1651), .B(n350), .Z(n188) );
  CND2XL U1773 ( .A(n430), .B(n415), .Z(n198) );
  CND2XL U1774 ( .A(n791), .B(n800), .Z(n334) );
  CND2IXL U1775 ( .B(n358), .A(n359), .Z(n190) );
  CND2IXL U1776 ( .B(n366), .A(n367), .Z(n192) );
  CND2XL U1777 ( .A(n1656), .B(n380), .Z(n195) );
  CND2XL U1778 ( .A(n1655), .B(n372), .Z(n193) );
  CND2XL U1779 ( .A(n1654), .B(n364), .Z(n191) );
  CEOXL U1780 ( .A(n376), .B(n194), .Z(product[3]) );
  CND2X1 U1781 ( .A(n662), .B(n649), .Z(n1676) );
  CENX1 U1782 ( .A(n1633), .B(n1667), .Z(n639) );
  CEOXL U1783 ( .A(n649), .B(n662), .Z(n1633) );
  CND2XL U1784 ( .A(n843), .B(n846), .Z(n367) );
  CEN3X1 U1785 ( .A(n434), .B(n1634), .C(n432), .Z(n415) );
  CEN3X2 U1786 ( .A(n436), .B(n418), .C(n417), .Z(n1634) );
  CAN2XL U1787 ( .A(n1566), .B(n383), .Z(product[1]) );
  CNR2IXL U1788 ( .B(n1687), .A(n58), .Z(n975) );
  COND2X1 U1789 ( .A(n53), .B(n1277), .C(n1276), .D(n50), .Z(n995) );
  CNR2IXL U1790 ( .B(n1687), .A(n89), .Z(n907) );
  CNR2IXL U1791 ( .B(n1687), .A(n1666), .Z(n921) );
  CNR2IXL U1792 ( .B(n1687), .A(n105), .Z(n877) );
  CNR2IXL U1793 ( .B(n1687), .A(n6), .Z(product[0]) );
  CENX4 U1794 ( .A(n1715), .B(a[12]), .Z(n58) );
  CENX4 U1795 ( .A(n1710), .B(a[10]), .Z(n50) );
  CND2X4 U1796 ( .A(n1458), .B(n6), .Z(n9) );
  CEOX2 U1797 ( .A(a[0]), .B(n1559), .Z(n1458) );
  CND2IX4 U1798 ( .B(n1635), .A(n24), .Z(n27) );
  CENX2 U1799 ( .A(n1721), .B(a[16]), .Z(n74) );
  CIVX4 U1800 ( .A(a[0]), .Z(n6) );
  CND2X2 U1801 ( .A(n1608), .B(n1446), .Z(n102) );
  CEOX1 U1802 ( .A(a[24]), .B(n1685), .Z(n1446) );
  CNIVX4 U1803 ( .A(n93), .Z(n1684) );
  CENX1 U1804 ( .A(a[8]), .B(n1712), .Z(n1637) );
  CND2XL U1805 ( .A(n1443), .B(n114), .Z(n115) );
  COND1XL U1806 ( .A(n223), .B(n1596), .C(n226), .Z(n222) );
  CAOR1X1 U1807 ( .A(n210), .B(n1641), .C(n205), .Z(n1638) );
  CANR1XL U1808 ( .A(n390), .B(n241), .C(n238), .Z(n236) );
  CANR1XL U1809 ( .A(n228), .B(n241), .C(n229), .Z(n227) );
  CNR2IXL U1810 ( .B(n228), .A(n223), .Z(n221) );
  COND1XL U1811 ( .A(n330), .B(n313), .C(n314), .Z(n312) );
  CND2X1 U1812 ( .A(n320), .B(n1645), .Z(n313) );
  CND2X1 U1813 ( .A(n1646), .B(n1644), .Z(n280) );
  CNR2X1 U1814 ( .A(n539), .B(n562), .Z(n234) );
  CANR1XL U1815 ( .A(n1647), .B(n264), .C(n257), .Z(n253) );
  CNR2X1 U1816 ( .A(n563), .B(n586), .Z(n239) );
  CENX1 U1817 ( .A(n297), .B(n179), .Z(product[18]) );
  CND2X1 U1818 ( .A(n397), .B(n296), .Z(n179) );
  CND2X1 U1819 ( .A(n1643), .B(n270), .Z(n175) );
  COND1XL U1820 ( .A(n272), .B(n278), .C(n273), .Z(n271) );
  CENX1 U1821 ( .A(n260), .B(n174), .Z(product[23]) );
  COND1XL U1822 ( .A(n261), .B(n278), .C(n262), .Z(n260) );
  CENX1 U1823 ( .A(n251), .B(n173), .Z(product[24]) );
  COND1XL U1824 ( .A(n252), .B(n278), .C(n253), .Z(n251) );
  CND2X1 U1825 ( .A(n263), .B(n1647), .Z(n252) );
  CENX1 U1826 ( .A(n304), .B(n180), .Z(product[17]) );
  CND2X1 U1827 ( .A(n1642), .B(n303), .Z(n180) );
  COND1XL U1828 ( .A(n305), .B(n1565), .C(n306), .Z(n304) );
  CENX1 U1829 ( .A(n291), .B(n178), .Z(product[19]) );
  CANR1XL U1830 ( .A(n1644), .B(n291), .C(n288), .Z(n286) );
  CND2XL U1831 ( .A(n1665), .B(n219), .Z(n169) );
  CND2X1 U1832 ( .A(n401), .B(n323), .Z(n183) );
  CANR1XL U1833 ( .A(n402), .B(n329), .C(n326), .Z(n324) );
  COR2X1 U1834 ( .A(n459), .B(n486), .Z(n1640) );
  CND2X1 U1835 ( .A(n459), .B(n486), .Z(n212) );
  COR2X1 U1836 ( .A(n431), .B(n458), .Z(n1641) );
  CND2X1 U1837 ( .A(n431), .B(n458), .Z(n207) );
  COND1XL U1838 ( .A(n337), .B(n333), .C(n334), .Z(n332) );
  CND2X1 U1839 ( .A(n1652), .B(n1651), .Z(n340) );
  CNR2X1 U1840 ( .A(n767), .B(n778), .Z(n322) );
  CENX1 U1841 ( .A(n189), .B(n357), .Z(product[8]) );
  CENX1 U1842 ( .A(n188), .B(n351), .Z(product[9]) );
  CENX1 U1843 ( .A(n335), .B(n185), .Z(product[12]) );
  CND2X1 U1844 ( .A(n403), .B(n334), .Z(n185) );
  COND1XL U1845 ( .A(n336), .B(n338), .C(n337), .Z(n335) );
  CENX1 U1846 ( .A(n329), .B(n184), .Z(product[13]) );
  CNR2X1 U1847 ( .A(n739), .B(n752), .Z(n305) );
  COR2X1 U1848 ( .A(n723), .B(n738), .Z(n1642) );
  CEOX1 U1849 ( .A(n346), .B(n187), .Z(product[10]) );
  CANR1XL U1850 ( .A(n1651), .B(n351), .C(n348), .Z(n346) );
  CEOX1 U1851 ( .A(n186), .B(n338), .Z(product[11]) );
  COR2X1 U1852 ( .A(n631), .B(n650), .Z(n1643) );
  COR2X1 U1853 ( .A(n689), .B(n706), .Z(n1644) );
  COR2X1 U1854 ( .A(n753), .B(n766), .Z(n1645) );
  CND2X1 U1855 ( .A(n651), .B(n670), .Z(n273) );
  CND2X1 U1856 ( .A(n739), .B(n752), .Z(n306) );
  COR2X1 U1857 ( .A(n671), .B(n688), .Z(n1646) );
  CND2X1 U1858 ( .A(n707), .B(n722), .Z(n296) );
  COR2X1 U1859 ( .A(n609), .B(n630), .Z(n1647) );
  CND2X1 U1860 ( .A(n689), .B(n706), .Z(n290) );
  CND2X1 U1861 ( .A(n631), .B(n650), .Z(n270) );
  CND2X1 U1862 ( .A(n587), .B(n608), .Z(n250) );
  CND2X1 U1863 ( .A(n671), .B(n688), .Z(n285) );
  CND2X1 U1864 ( .A(n753), .B(n766), .Z(n318) );
  CND2X1 U1865 ( .A(n723), .B(n738), .Z(n303) );
  COR2X1 U1866 ( .A(n587), .B(n608), .Z(n1648) );
  CANR1XL U1867 ( .A(n381), .B(n1656), .C(n378), .Z(n376) );
  COND1XL U1868 ( .A(n358), .B(n360), .C(n359), .Z(n357) );
  CENX1 U1869 ( .A(n1649), .B(n633), .Z(n631) );
  CENX1 U1870 ( .A(n635), .B(n652), .Z(n1649) );
  CNR2X1 U1871 ( .A(n801), .B(n810), .Z(n336) );
  CNR2X1 U1872 ( .A(n791), .B(n800), .Z(n333) );
  CNR2X1 U1873 ( .A(n779), .B(n790), .Z(n327) );
  COR2X1 U1874 ( .A(n827), .B(n832), .Z(n1650) );
  COR2X1 U1875 ( .A(n811), .B(n818), .Z(n1652) );
  CND2X1 U1876 ( .A(n779), .B(n790), .Z(n328) );
  CND2X1 U1877 ( .A(n801), .B(n810), .Z(n337) );
  CND2X1 U1878 ( .A(n827), .B(n832), .Z(n356) );
  CND2X1 U1879 ( .A(n811), .B(n818), .Z(n345) );
  CND2X1 U1880 ( .A(n819), .B(n826), .Z(n350) );
  COR2X1 U1881 ( .A(n430), .B(n415), .Z(n1653) );
  CENX1 U1882 ( .A(n191), .B(n365), .Z(product[6]) );
  CENX1 U1883 ( .A(n193), .B(n373), .Z(product[4]) );
  CND2X1 U1884 ( .A(n412), .B(n375), .Z(n194) );
  CENX1 U1885 ( .A(n195), .B(n381), .Z(product[2]) );
  CNR2X1 U1886 ( .A(n833), .B(n838), .Z(n358) );
  CNR2X1 U1887 ( .A(n843), .B(n846), .Z(n366) );
  CNR2X1 U1888 ( .A(n849), .B(n1104), .Z(n374) );
  CND2X1 U1889 ( .A(n833), .B(n838), .Z(n359) );
  CND2X1 U1890 ( .A(n847), .B(n848), .Z(n372) );
  CND2X1 U1891 ( .A(n839), .B(n842), .Z(n364) );
  CND2X1 U1892 ( .A(n1135), .B(n1105), .Z(n380) );
  COR2X1 U1893 ( .A(n839), .B(n842), .Z(n1654) );
  COR2X1 U1894 ( .A(n847), .B(n848), .Z(n1655) );
  COR2X1 U1895 ( .A(n1135), .B(n1105), .Z(n1656) );
  CENX1 U1896 ( .A(n1721), .B(n1679), .Z(n1230) );
  CENX1 U1897 ( .A(n1715), .B(n1680), .Z(n1273) );
  CENX1 U1898 ( .A(n1715), .B(n1679), .Z(n1274) );
  CENX1 U1899 ( .A(n1688), .B(n1722), .Z(n1233) );
  CENX1 U1900 ( .A(n1721), .B(n1680), .Z(n1229) );
  CENX1 U1901 ( .A(n1562), .B(n1680), .Z(n1418) );
  CENX1 U1902 ( .A(n1562), .B(n1688), .Z(n1422) );
  CENX1 U1903 ( .A(n1562), .B(n1677), .Z(n1421) );
  CENX1 U1904 ( .A(n1562), .B(n1679), .Z(n1419) );
  CENX1 U1905 ( .A(n1562), .B(n1678), .Z(n1420) );
  CENX1 U1906 ( .A(n1673), .B(n1678), .Z(n1275) );
  CIVX2 U1907 ( .A(n1720), .Z(n1719) );
  CENX1 U1908 ( .A(n1715), .B(n1689), .Z(n1277) );
  CENX1 U1909 ( .A(n1715), .B(n1677), .Z(n1276) );
  CENX1 U1910 ( .A(n1698), .B(n1689), .Z(n1358) );
  CNR2IX1 U1911 ( .B(n1687), .A(n95), .Z(n895) );
  CNIVX1 U1912 ( .A(n15), .Z(n1662) );
  CNR2IX1 U1913 ( .B(n1687), .A(n1662), .Z(n1105) );
  CENX1 U1914 ( .A(n1699), .B(n1679), .Z(n1355) );
  CENX1 U1915 ( .A(n1699), .B(n1678), .Z(n1356) );
  CENX1 U1916 ( .A(n1709), .B(n1680), .Z(n1298) );
  CENX1 U1917 ( .A(n1709), .B(n1679), .Z(n1299) );
  CENX1 U1918 ( .A(n1698), .B(n1680), .Z(n1354) );
  CENX1 U1919 ( .A(n1705), .B(n1678), .Z(n1327) );
  CENX1 U1920 ( .A(n1722), .B(n1678), .Z(n1231) );
  CENX1 U1921 ( .A(n1722), .B(n1677), .Z(n1232) );
  CENX1 U1922 ( .A(n1682), .B(n1680), .Z(n1193) );
  CENX1 U1923 ( .A(n1678), .B(n1682), .Z(n1195) );
  CENX1 U1924 ( .A(n1682), .B(n1679), .Z(n1194) );
  CNIVX2 U1925 ( .A(n15), .Z(n1661) );
  CENX1 U1926 ( .A(n1693), .B(n1678), .Z(n1387) );
  CENX1 U1927 ( .A(n1693), .B(n1677), .Z(n1388) );
  CENX1 U1928 ( .A(n1693), .B(n1680), .Z(n1385) );
  CENX1 U1929 ( .A(n1693), .B(n1679), .Z(n1386) );
  CENX1 U1930 ( .A(n1688), .B(n1685), .Z(n1158) );
  CENX1 U1931 ( .A(n1679), .B(n1684), .Z(n1166) );
  CENX1 U1932 ( .A(n1677), .B(n1685), .Z(n1157) );
  CENX1 U1933 ( .A(n1677), .B(n1684), .Z(n1168) );
  CENX1 U1934 ( .A(n1678), .B(n1684), .Z(n1167) );
  CENX1 U1935 ( .A(n1688), .B(n1684), .Z(n1169) );
  CENX1 U1936 ( .A(n1680), .B(n1684), .Z(n1165) );
  CENX1 U1937 ( .A(n1678), .B(n1685), .Z(n1156) );
  CENX1 U1938 ( .A(n1679), .B(n1685), .Z(n1155) );
  CENX1 U1939 ( .A(n1680), .B(n1685), .Z(n1154) );
  CENX1 U1940 ( .A(n1688), .B(n1682), .Z(n1197) );
  CENX1 U1941 ( .A(n1705), .B(n1679), .Z(n1326) );
  CENX1 U1942 ( .A(n1705), .B(n1680), .Z(n1325) );
  CENX1 U1943 ( .A(n1705), .B(n1677), .Z(n1328) );
  CENX1 U1944 ( .A(n1686), .B(n1705), .Z(n1330) );
  CENX1 U1945 ( .A(n1686), .B(n1682), .Z(n1198) );
  CENX1 U1946 ( .A(n1686), .B(n1712), .Z(n1303) );
  CENX1 U1947 ( .A(n1705), .B(n1688), .Z(n1329) );
  CNR2IX1 U1948 ( .B(n1687), .A(n24), .Z(n1075) );
  COND2X1 U1949 ( .A(n27), .B(n1348), .C(n1347), .D(n24), .Z(n1063) );
  CNR2IX1 U1950 ( .B(n1687), .A(n42), .Z(n1021) );
  CNR2IX1 U1951 ( .B(n1687), .A(n33), .Z(n1047) );
  COND2X1 U1952 ( .A(n27), .B(n1358), .C(n1357), .D(n24), .Z(n1073) );
  CEOX1 U1953 ( .A(n872), .B(n886), .Z(n429) );
  CENX1 U1954 ( .A(n1707), .B(n153), .Z(n1311) );
  CENX1 U1955 ( .A(n1682), .B(n132), .Z(n1191) );
  CENX1 U1956 ( .A(n1722), .B(n138), .Z(n1224) );
  CENX1 U1957 ( .A(n1707), .B(n152), .Z(n1312) );
  CENX1 U1958 ( .A(n1705), .B(n151), .Z(n1313) );
  CENX1 U1959 ( .A(n1701), .B(n151), .Z(n1342) );
  CENX1 U1960 ( .A(n1701), .B(n152), .Z(n1341) );
  CENX1 U1961 ( .A(n1711), .B(n136), .Z(n1294) );
  CENX1 U1962 ( .A(n1682), .B(n136), .Z(n1189) );
  CENX1 U1963 ( .A(n1723), .B(n146), .Z(n1220) );
  CENX1 U1964 ( .A(n1682), .B(n142), .Z(n1186) );
  CENX1 U1965 ( .A(n1723), .B(n148), .Z(n1219) );
  CENX1 U1966 ( .A(n1711), .B(n151), .Z(n1286) );
  CENX1 U1967 ( .A(n1682), .B(n138), .Z(n1188) );
  CENX1 U1968 ( .A(n1695), .B(n152), .Z(n1372) );
  CENX1 U1969 ( .A(n1694), .B(n151), .Z(n1373) );
  CENX1 U1970 ( .A(n1562), .B(n152), .Z(n1405) );
  CENX1 U1971 ( .A(n1693), .B(n156), .Z(n1368) );
  CENX1 U1972 ( .A(n1693), .B(n157), .Z(n1367) );
  CENX1 U1973 ( .A(n1696), .B(n142), .Z(n1378) );
  CENX1 U1974 ( .A(n1694), .B(b[24]), .Z(n1366) );
  CENX1 U1975 ( .A(n1692), .B(b[26]), .Z(n1364) );
  CENX1 U1976 ( .A(n1692), .B(b[27]), .Z(n1363) );
  CENX1 U1977 ( .A(n1692), .B(b[28]), .Z(n1362) );
  CENX1 U1978 ( .A(n104), .B(a[28]), .Z(n110) );
  CENX1 U1979 ( .A(n1699), .B(b[27]), .Z(n1332) );
  CENX1 U1980 ( .A(n1562), .B(b[31]), .Z(n1392) );
  CENX1 U1981 ( .A(n1678), .B(n109), .Z(n1140) );
  CENX1 U1982 ( .A(n109), .B(a[30]), .Z(n114) );
  CENX1 U1983 ( .A(n1709), .B(n157), .Z(n1280) );
  CENX1 U1984 ( .A(n1707), .B(n146), .Z(n1316) );
  CENX1 U1985 ( .A(n1699), .B(n155), .Z(n1338) );
  CENX1 U1986 ( .A(n1699), .B(n154), .Z(n1339) );
  CENX1 U1987 ( .A(n1707), .B(n148), .Z(n1315) );
  CENX1 U1988 ( .A(n1699), .B(n157), .Z(n1336) );
  CENX1 U1989 ( .A(n1699), .B(n156), .Z(n1337) );
  CENX1 U1990 ( .A(n1704), .B(n154), .Z(n1310) );
  CENX1 U1991 ( .A(n1709), .B(n154), .Z(n1283) );
  CENX1 U1992 ( .A(n1711), .B(n155), .Z(n1282) );
  CENX1 U1993 ( .A(n1709), .B(n153), .Z(n1284) );
  CENX1 U1994 ( .A(n1698), .B(b[24]), .Z(n1335) );
  CENX1 U1995 ( .A(n1709), .B(n156), .Z(n1281) );
  CENX1 U1996 ( .A(n1698), .B(b[26]), .Z(n1333) );
  CENX1 U1997 ( .A(n1696), .B(n146), .Z(n1376) );
  CENX1 U1998 ( .A(n1677), .B(n104), .Z(n1148) );
  CENX1 U1999 ( .A(n1679), .B(n104), .Z(n1146) );
  CENX1 U2000 ( .A(n1678), .B(n104), .Z(n1147) );
  CENX1 U2001 ( .A(n1693), .B(n155), .Z(n1369) );
  CENX1 U2002 ( .A(n1693), .B(n154), .Z(n1370) );
  CENX1 U2003 ( .A(n1696), .B(n148), .Z(n1375) );
  CENX1 U2004 ( .A(n1688), .B(n104), .Z(n1149) );
  CENX1 U2005 ( .A(n1704), .B(n155), .Z(n1309) );
  CENX1 U2006 ( .A(n1680), .B(n104), .Z(n1145) );
  CENX1 U2007 ( .A(n1686), .B(n113), .Z(n1138) );
  CENX1 U2008 ( .A(n1688), .B(n113), .Z(n1137) );
  CENX1 U2009 ( .A(n1686), .B(n104), .Z(n1150) );
  CENX1 U2010 ( .A(n1686), .B(n109), .Z(n1143) );
  CIVX2 U2011 ( .A(n63), .Z(n1724) );
  CENX1 U2012 ( .A(n1681), .B(a[18]), .Z(n82) );
  CIVX2 U2013 ( .A(n39), .Z(n1713) );
  CND2X1 U2014 ( .A(n1444), .B(n110), .Z(n112) );
  CEOXL U2015 ( .A(a[28]), .B(n109), .Z(n1444) );
  CNIVX4 U2016 ( .A(n99), .Z(n1685) );
  CEOX1 U2017 ( .A(a[30]), .B(n113), .Z(n1443) );
  CENX1 U2018 ( .A(n1691), .B(a[2]), .Z(n15) );
  CAN2XL U2019 ( .A(n1641), .B(n207), .Z(n1663) );
  CENX1 U2020 ( .A(n1698), .B(n1677), .Z(n1357) );
  COND2XL U2021 ( .A(n53), .B(n1258), .C(n1257), .D(n50), .Z(n976) );
  CNR2IXL U2022 ( .B(n1687), .A(n50), .Z(n997) );
  COND2XL U2023 ( .A(n53), .B(n1261), .C(n1260), .D(n50), .Z(n979) );
  COND2XL U2024 ( .A(n53), .B(n1269), .C(n1268), .D(n50), .Z(n987) );
  COND2XL U2025 ( .A(n53), .B(n1260), .C(n1259), .D(n50), .Z(n978) );
  COND2XL U2026 ( .A(n1278), .B(n53), .C(n1277), .D(n50), .Z(n996) );
  COND2XL U2027 ( .A(n53), .B(n1271), .C(n1270), .D(n50), .Z(n989) );
  COND2XL U2028 ( .A(n53), .B(n1270), .C(n1269), .D(n50), .Z(n988) );
  CANR1XL U2029 ( .A(n320), .B(n329), .C(n321), .Z(n319) );
  COND2XL U2030 ( .A(n61), .B(n1720), .C(n58), .D(n1256), .Z(n859) );
  CIVXL U2031 ( .A(n1691), .Z(n1664) );
  COR2XL U2032 ( .A(n512), .B(n487), .Z(n1665) );
  CIVXL U2033 ( .A(n647), .Z(n1667) );
  CND2XL U2034 ( .A(n1647), .B(n259), .Z(n174) );
  CIVX1 U2035 ( .A(n259), .Z(n257) );
  COND2X1 U2036 ( .A(n77), .B(n1212), .C(n1211), .D(n1619), .Z(n933) );
  CND2XL U2037 ( .A(n633), .B(n652), .Z(n1670) );
  CND2X1 U2038 ( .A(n633), .B(n635), .Z(n1671) );
  CND2XL U2039 ( .A(n652), .B(n635), .Z(n1672) );
  CND3XL U2040 ( .A(n1670), .B(n1671), .C(n1672), .Z(n630) );
  CND2X1 U2041 ( .A(n609), .B(n630), .Z(n259) );
  CENX1 U2042 ( .A(n1698), .B(n142), .Z(n1347) );
  CENX1 U2043 ( .A(n1706), .B(n142), .Z(n1318) );
  CENX1 U2044 ( .A(n1711), .B(n142), .Z(n1291) );
  CIVX1 U2045 ( .A(n1713), .Z(n1709) );
  CNIVX1 U2046 ( .A(n120), .Z(n1689) );
  CND2X1 U2047 ( .A(n647), .B(n662), .Z(n1674) );
  COND2X1 U2048 ( .A(n27), .B(n1342), .C(n1341), .D(n24), .Z(n1057) );
  CIVX1 U2049 ( .A(n1714), .Z(n1712) );
  COND2XL U2050 ( .A(n9), .B(n1664), .C(n6), .D(n1424), .Z(n865) );
  CND2IXL U2051 ( .B(n1687), .A(n1560), .Z(n1424) );
  CND2X1 U2052 ( .A(n1136), .B(n865), .Z(n383) );
  COND2X1 U2053 ( .A(n77), .B(n1207), .C(n1206), .D(n1619), .Z(n928) );
  COND2X1 U2054 ( .A(n77), .B(n1214), .C(n1213), .D(n1619), .Z(n935) );
  COND2X1 U2055 ( .A(n77), .B(n1206), .C(n1205), .D(n1619), .Z(n927) );
  COND2X1 U2056 ( .A(n77), .B(n1205), .C(n1204), .D(n1619), .Z(n926) );
  CFA1XL U2057 ( .A(n1036), .B(n737), .CI(n1062), .CO(n730), .S(n731) );
  CND2X1 U2058 ( .A(n647), .B(n649), .Z(n1675) );
  COND2XL U2059 ( .A(n53), .B(n1717), .C(n50), .D(n1279), .Z(n860) );
  COND1XL U2060 ( .A(n298), .B(n1565), .C(n299), .Z(n297) );
  COND2XL U2061 ( .A(n27), .B(n1703), .C(n24), .D(n1360), .Z(n863) );
  COND2X1 U2062 ( .A(n1668), .B(n1328), .C(n1327), .D(n33), .Z(n1044) );
  CIVX1 U2063 ( .A(n1708), .Z(n1705) );
  COND2X1 U2064 ( .A(n77), .B(n1211), .C(n1210), .D(n1619), .Z(n932) );
  CIVX1 U2065 ( .A(n1703), .Z(n1700) );
  COND2XL U2066 ( .A(n18), .B(n1697), .C(n1661), .D(n1391), .Z(n864) );
  CIVX1 U2067 ( .A(n1697), .Z(n1696) );
  CIVX1 U2068 ( .A(n1708), .Z(n1707) );
  CND2IXL U2069 ( .B(n1687), .A(n1692), .Z(n1391) );
  CENX1 U2070 ( .A(n1705), .B(n156), .Z(n1308) );
  CND2IXL U2071 ( .B(n1687), .A(n1707), .Z(n1331) );
  CENX1 U2072 ( .A(n1707), .B(n157), .Z(n1307) );
  CENX1 U2073 ( .A(n1705), .B(b[24]), .Z(n1306) );
  COND2X1 U2074 ( .A(n69), .B(n1226), .C(n1225), .D(n66), .Z(n946) );
  COND2XL U2075 ( .A(n1668), .B(n1306), .C(n1305), .D(n33), .Z(n1022) );
  COND2XL U2076 ( .A(n1668), .B(n1308), .C(n1307), .D(n33), .Z(n1024) );
  COND2XL U2077 ( .A(n1669), .B(n1307), .C(n1306), .D(n33), .Z(n1023) );
  COND2XL U2078 ( .A(n1668), .B(n1322), .C(n1321), .D(n33), .Z(n1038) );
  COND2XL U2079 ( .A(n1668), .B(n1326), .C(n1325), .D(n33), .Z(n1042) );
  COND2XL U2080 ( .A(n1668), .B(n1708), .C(n33), .D(n1331), .Z(n862) );
  COND2XL U2081 ( .A(n1330), .B(n1669), .C(n1329), .D(n33), .Z(n1046) );
  COND2XL U2082 ( .A(n1668), .B(n1320), .C(n1319), .D(n33), .Z(n1036) );
  CENX1 U2083 ( .A(n1711), .B(n146), .Z(n1289) );
  CENX1 U2084 ( .A(n1711), .B(n148), .Z(n1288) );
  CIVX2 U2085 ( .A(n1724), .Z(n1722) );
  CIVX1 U2086 ( .A(n1703), .Z(n1699) );
  CND2XL U2087 ( .A(n216), .B(n228), .Z(n214) );
  CEOXL U2088 ( .A(n360), .B(n190), .Z(product[7]) );
  CEOXL U2089 ( .A(n368), .B(n192), .Z(product[5]) );
  CIVX1 U2090 ( .A(n1703), .Z(n1698) );
  COND2X1 U2091 ( .A(n77), .B(n1210), .C(n1209), .D(n1619), .Z(n931) );
  COND2XL U2092 ( .A(n77), .B(n1201), .C(n1200), .D(n1619), .Z(n922) );
  COND2XL U2093 ( .A(n77), .B(n1204), .C(n1203), .D(n1619), .Z(n925) );
  COND2XL U2094 ( .A(n1215), .B(n77), .C(n1619), .D(n1214), .Z(n936) );
  COND2XL U2095 ( .A(n77), .B(n1203), .C(n1202), .D(n1619), .Z(n924) );
  COND2XL U2096 ( .A(n77), .B(n1202), .C(n1201), .D(n1619), .Z(n923) );
  COND2XL U2097 ( .A(n77), .B(n1213), .C(n1212), .D(n1619), .Z(n934) );
  COND2XL U2098 ( .A(n77), .B(n1475), .C(n1619), .D(n1216), .Z(n857) );
  CND2IXL U2099 ( .B(n1687), .A(n1721), .Z(n1235) );
  CND2X4 U2100 ( .A(n1457), .B(n1660), .Z(n18) );
  CIVXL U2101 ( .A(n1697), .Z(n1692) );
  CIVXL U2102 ( .A(n1697), .Z(n1695) );
  CIVXL U2103 ( .A(n1703), .Z(n1701) );
  CIVXL U2104 ( .A(n1708), .Z(n1706) );
  CIVXL U2105 ( .A(n1724), .Z(n1723) );
  CIVX2 U2106 ( .A(n374), .Z(n412) );
  CIVX2 U2107 ( .A(n336), .Z(n404) );
  CIVX2 U2108 ( .A(n333), .Z(n403) );
  CIVX2 U2109 ( .A(n295), .Z(n397) );
  CIVX2 U2110 ( .A(n383), .Z(n381) );
  CIVX2 U2111 ( .A(n380), .Z(n378) );
  CIVX2 U2112 ( .A(n372), .Z(n370) );
  CIVX2 U2113 ( .A(n364), .Z(n362) );
  CIVX2 U2114 ( .A(n356), .Z(n354) );
  CIVX2 U2115 ( .A(n350), .Z(n348) );
  CIVX2 U2116 ( .A(n345), .Z(n343) );
  CIVX2 U2117 ( .A(n339), .Z(n338) );
  CIVX2 U2118 ( .A(n328), .Z(n326) );
  CIVX2 U2119 ( .A(n327), .Z(n402) );
  CIVX2 U2120 ( .A(n318), .Z(n316) );
  CIVX2 U2121 ( .A(n306), .Z(n308) );
  CIVX2 U2122 ( .A(n305), .Z(n399) );
  CIVX2 U2123 ( .A(n290), .Z(n288) );
  CIVX2 U2124 ( .A(n285), .Z(n283) );
  CIVX2 U2125 ( .A(n272), .Z(n394) );
  CIVX2 U2126 ( .A(n270), .Z(n268) );
  CIVX2 U2127 ( .A(n261), .Z(n263) );
  CIVX2 U2128 ( .A(n250), .Z(n248) );
  CIVX2 U2129 ( .A(n240), .Z(n238) );
  CIVX2 U2130 ( .A(n239), .Z(n390) );
  CIVX2 U2131 ( .A(n212), .Z(n210) );
  CIVX2 U2132 ( .A(n207), .Z(n205) );
  CIVX2 U2133 ( .A(n1681), .Z(n1475) );
  CIVX2 U2134 ( .A(n104), .Z(n1470) );
  CIVX2 U2135 ( .A(n109), .Z(n1469) );
  CIVX2 U2136 ( .A(n113), .Z(n1468) );
endmodule


module calc_DW_mult_uns_17 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n3, n9, n12, n18, n21, n27, n30, n33, n36, n39, n42, n44, n48, n50,
         n53, n55, n58, n61, n63, n66, n69, n71, n74, n77, n79, n82, n85, n87,
         n89, n91, n93, n95, n97, n99, n100, n102, n104, n105, n107, n109,
         n110, n112, n113, n114, n115, n116, n120, n122, n124, n126, n128,
         n130, n132, n134, n136, n138, n140, n142, n144, n146, n148, n150,
         n151, n152, n153, n154, n155, n156, n157, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n198, n199, n206, n207, n210, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n226, n227,
         n228, n229, n231, n234, n235, n236, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n249, n250, n251, n252, n253, n257, n259,
         n260, n261, n262, n263, n264, n268, n270, n271, n272, n273, n275,
         n278, n279, n280, n281, n283, n285, n286, n288, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n301, n303, n304, n305,
         n306, n308, n312, n313, n314, n316, n318, n319, n320, n321, n322,
         n323, n324, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n343, n345, n346, n348,
         n350, n351, n352, n354, n356, n357, n358, n359, n360, n362, n364,
         n365, n366, n367, n368, n370, n372, n373, n374, n375, n376, n378,
         n380, n381, n383, n385, n387, n388, n390, n391, n394, n397, n399,
         n401, n402, n403, n404, n412, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1443, n1445, n1446, n1447, n1448, n1449, n1451, n1452, n1454,
         n1455, n1456, n1458, n1468, n1469, n1470, n1473, n1474, n1475, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736;
  assign n3 = a[1];
  assign n12 = a[3];
  assign n21 = a[5];
  assign n30 = a[7];
  assign n39 = a[9];
  assign n48 = a[11];
  assign n55 = a[13];
  assign n63 = a[15];
  assign n71 = a[17];
  assign n79 = a[19];
  assign n87 = a[21];
  assign n93 = a[23];
  assign n99 = a[25];
  assign n104 = a[27];
  assign n109 = a[29];
  assign n113 = a[31];
  assign n116 = b[0];
  assign n120 = b[1];
  assign n122 = b[2];
  assign n124 = b[3];
  assign n126 = b[4];
  assign n128 = b[5];
  assign n130 = b[6];
  assign n132 = b[7];
  assign n134 = b[8];
  assign n136 = b[9];
  assign n138 = b[10];
  assign n140 = b[11];
  assign n142 = b[12];
  assign n144 = b[13];
  assign n146 = b[14];
  assign n148 = b[15];
  assign n150 = b[16];
  assign n151 = b[17];
  assign n152 = b[18];
  assign n153 = b[19];
  assign n154 = b[20];
  assign n155 = b[21];
  assign n156 = b[22];
  assign n157 = b[23];

  CNR2X2 U171 ( .A(n513), .B(n538), .Z(n223) );
  CND2X2 U192 ( .A(n563), .B(n586), .Z(n240) );
  CNR2X2 U204 ( .A(n587), .B(n608), .Z(n249) );
  CND2X2 U241 ( .A(n651), .B(n670), .Z(n273) );
  CEO3X2 U412 ( .A(n444), .B(n423), .C(n442), .Z(n419) );
  CEO3X2 U413 ( .A(n425), .B(n424), .C(n446), .Z(n420) );
  CEO3X2 U414 ( .A(n428), .B(n427), .C(n426), .Z(n421) );
  CEO3X2 U416 ( .A(n456), .B(n429), .C(n454), .Z(n423) );
  CEO3X2 U417 ( .A(n998), .B(n1022), .C(n1106), .Z(n424) );
  CEO3X2 U418 ( .A(n866), .B(n976), .C(n1076), .Z(n425) );
  CEO3X2 U419 ( .A(n922), .B(n938), .C(n1048), .Z(n426) );
  CEO3X2 U420 ( .A(n850), .B(n896), .C(n956), .Z(n427) );
  CEO3X2 U421 ( .A(n878), .B(n868), .C(n908), .Z(n428) );
  CFA1X1 U423 ( .A(n435), .B(n433), .CI(n460), .CO(n430), .S(n431) );
  CFA1X1 U424 ( .A(n439), .B(n462), .CI(n437), .CO(n432), .S(n433) );
  CFA1X1 U425 ( .A(n441), .B(n464), .CI(n466), .CO(n434), .S(n435) );
  CFA1X1 U426 ( .A(n445), .B(n443), .CI(n468), .CO(n436), .S(n437) );
  CFA1X1 U427 ( .A(n472), .B(n447), .CI(n470), .CO(n438), .S(n439) );
  CFA1X1 U428 ( .A(n474), .B(n449), .CI(n451), .CO(n440), .S(n441) );
  CFA1X1 U429 ( .A(n457), .B(n453), .CI(n455), .CO(n442), .S(n443) );
  CFA1X1 U430 ( .A(n480), .B(n476), .CI(n478), .CO(n444), .S(n445) );
  CFA1X1 U431 ( .A(n1023), .B(n482), .CI(n484), .CO(n446), .S(n447) );
  CFA1X1 U432 ( .A(n957), .B(n1077), .CI(n1107), .CO(n448), .S(n449) );
  CFA1X1 U433 ( .A(n939), .B(n1049), .CI(n999), .CO(n450), .S(n451) );
  CFA1X1 U435 ( .A(n869), .B(n909), .CI(n887), .CO(n454), .S(n455) );
  CFA1X1 U436 ( .A(n867), .B(n879), .CI(n873), .CO(n456), .S(n457) );
  CFA1X1 U437 ( .A(n463), .B(n461), .CI(n488), .CO(n458), .S(n459) );
  CFA1X1 U438 ( .A(n467), .B(n490), .CI(n465), .CO(n460), .S(n461) );
  CFA1X1 U439 ( .A(n469), .B(n492), .CI(n494), .CO(n462), .S(n463) );
  CFA1X1 U440 ( .A(n473), .B(n471), .CI(n496), .CO(n464), .S(n465) );
  CFA1X1 U441 ( .A(n475), .B(n498), .CI(n500), .CO(n466), .S(n467) );
  CFA1X1 U442 ( .A(n481), .B(n477), .CI(n479), .CO(n468), .S(n469) );
  CFA1X1 U443 ( .A(n502), .B(n483), .CI(n504), .CO(n470), .S(n471) );
  CFA1X1 U444 ( .A(n510), .B(n506), .CI(n508), .CO(n472), .S(n473) );
  CFA1X1 U445 ( .A(n1024), .B(n485), .CI(n1108), .CO(n474), .S(n475) );
  CFA1X1 U446 ( .A(n940), .B(n1050), .CI(n1000), .CO(n476), .S(n477) );
  CFA1X1 U447 ( .A(n870), .B(n1078), .CI(n958), .CO(n478), .S(n479) );
  CFA1X1 U448 ( .A(n898), .B(n978), .CI(n924), .CO(n480), .S(n481) );
  CHA1X1 U450 ( .A(n874), .B(n888), .CO(n484), .S(n485) );
  CFA1X1 U451 ( .A(n491), .B(n489), .CI(n514), .CO(n486), .S(n487) );
  CFA1X1 U452 ( .A(n495), .B(n516), .CI(n493), .CO(n488), .S(n489) );
  CFA1X1 U453 ( .A(n497), .B(n518), .CI(n520), .CO(n490), .S(n491) );
  CFA1X1 U454 ( .A(n501), .B(n499), .CI(n522), .CO(n492), .S(n493) );
  CFA1X1 U455 ( .A(n503), .B(n524), .CI(n526), .CO(n494), .S(n495) );
  CFA1X1 U456 ( .A(n509), .B(n505), .CI(n507), .CO(n496), .S(n497) );
  CFA1X1 U457 ( .A(n530), .B(n511), .CI(n528), .CO(n498), .S(n499) );
  CFA1X1 U458 ( .A(n536), .B(n532), .CI(n534), .CO(n500), .S(n501) );
  CFA1X1 U459 ( .A(n979), .B(n1079), .CI(n1001), .CO(n502), .S(n503) );
  CFA1X1 U460 ( .A(n959), .B(n1051), .CI(n1109), .CO(n504), .S(n505) );
  CFA1X1 U463 ( .A(n871), .B(n875), .CI(n881), .CO(n510), .S(n511) );
  CFA1X1 U464 ( .A(n517), .B(n515), .CI(n540), .CO(n512), .S(n513) );
  CFA1X1 U465 ( .A(n521), .B(n542), .CI(n519), .CO(n514), .S(n515) );
  CFA1X1 U466 ( .A(n546), .B(n544), .CI(n523), .CO(n516), .S(n517) );
  CFA1X1 U467 ( .A(n527), .B(n525), .CI(n548), .CO(n518), .S(n519) );
  CFA1X1 U468 ( .A(n533), .B(n550), .CI(n529), .CO(n520), .S(n521) );
  CFA1X1 U469 ( .A(n535), .B(n531), .CI(n552), .CO(n522), .S(n523) );
  CFA1X1 U470 ( .A(n558), .B(n554), .CI(n556), .CO(n524), .S(n525) );
  CFA1X1 U471 ( .A(n1002), .B(n560), .CI(n537), .CO(n526), .S(n527) );
  CFA1X1 U473 ( .A(n926), .B(n1052), .CI(n1619), .CO(n530), .S(n531) );
  CFA1X1 U474 ( .A(n1621), .B(n1026), .CI(n876), .CO(n532), .S(n533) );
  CFA1X1 U475 ( .A(n890), .B(n942), .CI(n900), .CO(n534), .S(n535) );
  CFA1X1 U477 ( .A(n543), .B(n541), .CI(n564), .CO(n538), .S(n539) );
  CFA1X1 U478 ( .A(n568), .B(n566), .CI(n545), .CO(n540), .S(n541) );
  CFA1X1 U479 ( .A(n570), .B(n547), .CI(n549), .CO(n542), .S(n543) );
  CFA1X1 U481 ( .A(n557), .B(n553), .CI(n555), .CO(n546), .S(n547) );
  CFA1X1 U482 ( .A(n578), .B(n559), .CI(n561), .CO(n548), .S(n549) );
  CFA1X1 U483 ( .A(n582), .B(n576), .CI(n580), .CO(n550), .S(n551) );
  CFA1X1 U484 ( .A(n1003), .B(n584), .CI(n1081), .CO(n552), .S(n553) );
  CFA1X1 U485 ( .A(n1053), .B(n961), .CI(n1111), .CO(n554), .S(n555) );
  CFA1X1 U486 ( .A(n913), .B(n1027), .CI(n943), .CO(n556), .S(n557) );
  CFA1X1 U487 ( .A(n901), .B(n981), .CI(n927), .CO(n558), .S(n559) );
  CFA1X1 U488 ( .A(n877), .B(n891), .CI(n883), .CO(n560), .S(n561) );
  CFA1X1 U489 ( .A(n567), .B(n565), .CI(n588), .CO(n562), .S(n563) );
  CFA1X1 U490 ( .A(n592), .B(n590), .CI(n569), .CO(n564), .S(n565) );
  CFA1X1 U491 ( .A(n594), .B(n571), .CI(n573), .CO(n566), .S(n567) );
  CFA1X1 U492 ( .A(n598), .B(n575), .CI(n596), .CO(n568), .S(n569) );
  CFA1X1 U493 ( .A(n581), .B(n577), .CI(n579), .CO(n570), .S(n571) );
  CFA1X1 U495 ( .A(n585), .B(n604), .CI(n606), .CO(n574), .S(n575) );
  CFA1X1 U499 ( .A(n853), .B(n962), .CI(n914), .CO(n582), .S(n583) );
  CHA1X1 U500 ( .A(n902), .B(n892), .CO(n584), .S(n585) );
  CFA1X1 U502 ( .A(n614), .B(n612), .CI(n593), .CO(n588), .S(n589) );
  CFA1X1 U503 ( .A(n616), .B(n595), .CI(n597), .CO(n590), .S(n591) );
  CFA1X1 U504 ( .A(n620), .B(n599), .CI(n618), .CO(n592), .S(n593) );
  CFA1X1 U505 ( .A(n605), .B(n601), .CI(n603), .CO(n594), .S(n595) );
  CFA1X1 U506 ( .A(n624), .B(n607), .CI(n622), .CO(n596), .S(n597) );
  CFA1X1 U507 ( .A(n1005), .B(n626), .CI(n628), .CO(n598), .S(n599) );
  CFA1X1 U508 ( .A(n983), .B(n1055), .CI(n1113), .CO(n600), .S(n601) );
  CFA1X1 U510 ( .A(n915), .B(n1029), .CI(n945), .CO(n604), .S(n605) );
  CFA1X1 U511 ( .A(n885), .B(n903), .CI(n893), .CO(n606), .S(n607) );
  CFA1X1 U512 ( .A(n613), .B(n611), .CI(n632), .CO(n608), .S(n609) );
  CFA1X1 U513 ( .A(n617), .B(n634), .CI(n615), .CO(n610), .S(n611) );
  CFA1X1 U514 ( .A(n638), .B(n636), .CI(n619), .CO(n612), .S(n613) );
  CFA1X1 U515 ( .A(n623), .B(n640), .CI(n621), .CO(n614), .S(n615) );
  CFA1X1 U516 ( .A(n642), .B(n625), .CI(n627), .CO(n616), .S(n617) );
  CFA1X1 U517 ( .A(n648), .B(n644), .CI(n646), .CO(n618), .S(n619) );
  CFA1X1 U520 ( .A(n894), .B(n1084), .CI(n964), .CO(n624), .S(n625) );
  CHA1X1 U522 ( .A(n854), .B(n916), .CO(n628), .S(n629) );
  CFA1X1 U524 ( .A(n639), .B(n654), .CI(n637), .CO(n632), .S(n633) );
  CFA1X1 U525 ( .A(n658), .B(n656), .CI(n641), .CO(n634), .S(n635) );
  CFA1X1 U526 ( .A(n645), .B(n660), .CI(n643), .CO(n636), .S(n637) );
  CFA1X1 U527 ( .A(n662), .B(n647), .CI(n649), .CO(n638), .S(n639) );
  CFA1X1 U528 ( .A(n668), .B(n664), .CI(n666), .CO(n640), .S(n641) );
  CFA1X1 U529 ( .A(n985), .B(n1115), .CI(n1031), .CO(n642), .S(n643) );
  CFA1X1 U530 ( .A(n947), .B(n1085), .CI(n1007), .CO(n644), .S(n645) );
  CFA1X1 U531 ( .A(n931), .B(n1617), .CI(n1678), .CO(n646), .S(n647) );
  CFA1X1 U532 ( .A(n895), .B(n917), .CI(n905), .CO(n648), .S(n649) );
  CFA1X1 U533 ( .A(n655), .B(n653), .CI(n672), .CO(n650), .S(n651) );
  CFA1X1 U534 ( .A(n659), .B(n674), .CI(n657), .CO(n652), .S(n653) );
  CFA1X1 U535 ( .A(n678), .B(n676), .CI(n661), .CO(n654), .S(n655) );
  CFA1X1 U536 ( .A(n680), .B(n663), .CI(n665), .CO(n656), .S(n657) );
  CFA1X1 U537 ( .A(n684), .B(n667), .CI(n682), .CO(n658), .S(n659) );
  CFA1X1 U538 ( .A(n1008), .B(n686), .CI(n669), .CO(n660), .S(n661) );
  CFA1X1 U541 ( .A(n918), .B(n1032), .CI(n948), .CO(n666), .S(n667) );
  CHA1X1 U542 ( .A(n855), .B(n932), .CO(n668), .S(n669) );
  CFA1X1 U543 ( .A(n675), .B(n673), .CI(n690), .CO(n670), .S(n671) );
  CFA1X1 U544 ( .A(n679), .B(n692), .CI(n677), .CO(n672), .S(n673) );
  CFA1X1 U545 ( .A(n681), .B(n694), .CI(n696), .CO(n674), .S(n675) );
  CFA1X1 U546 ( .A(n687), .B(n683), .CI(n685), .CO(n676), .S(n677) );
  CFA1X1 U547 ( .A(n702), .B(n698), .CI(n700), .CO(n678), .S(n679) );
  CFA1X1 U548 ( .A(n987), .B(n704), .CI(n1033), .CO(n680), .S(n681) );
  CFA1X1 U550 ( .A(n949), .B(n1615), .CI(n1009), .CO(n684), .S(n685) );
  CFA1X1 U551 ( .A(n907), .B(n933), .CI(n919), .CO(n686), .S(n687) );
  CFA1X1 U552 ( .A(n693), .B(n691), .CI(n708), .CO(n688), .S(n689) );
  CFA1X1 U553 ( .A(n697), .B(n710), .CI(n695), .CO(n690), .S(n691) );
  CFA1X1 U554 ( .A(n699), .B(n712), .CI(n714), .CO(n692), .S(n693) );
  CFA1X1 U555 ( .A(n718), .B(n701), .CI(n703), .CO(n694), .S(n695) );
  CFA1X1 U556 ( .A(n705), .B(n716), .CI(n720), .CO(n696), .S(n697) );
  CFA1X1 U557 ( .A(n1010), .B(n1118), .CI(n1034), .CO(n698), .S(n699) );
  CFA1X1 U558 ( .A(n920), .B(n1088), .CI(n988), .CO(n700), .S(n701) );
  CFA1X1 U559 ( .A(n934), .B(n1060), .CI(n968), .CO(n702), .S(n703) );
  CHA1X1 U560 ( .A(n856), .B(n950), .CO(n704), .S(n705) );
  CFA1X1 U561 ( .A(n711), .B(n709), .CI(n724), .CO(n706), .S(n707) );
  CFA1X1 U562 ( .A(n715), .B(n726), .CI(n713), .CO(n708), .S(n709) );
  CFA1X1 U563 ( .A(n717), .B(n728), .CI(n730), .CO(n710), .S(n711) );
  CFA1X1 U564 ( .A(n732), .B(n719), .CI(n721), .CO(n712), .S(n713) );
  CFA1X1 U565 ( .A(n1011), .B(n734), .CI(n736), .CO(n714), .S(n715) );
  CFA1X1 U566 ( .A(n989), .B(n1035), .CI(n1089), .CO(n716), .S(n717) );
  CFA1X1 U568 ( .A(n921), .B(n951), .CI(n935), .CO(n720), .S(n721) );
  CFA1X1 U569 ( .A(n727), .B(n725), .CI(n740), .CO(n722), .S(n723) );
  CFA1X1 U570 ( .A(n744), .B(n742), .CI(n729), .CO(n724), .S(n725) );
  CFA1X1 U571 ( .A(n735), .B(n731), .CI(n733), .CO(n726), .S(n727) );
  CFA1X1 U572 ( .A(n750), .B(n748), .CI(n746), .CO(n728), .S(n729) );
  CFA1X1 U573 ( .A(n970), .B(n737), .CI(n1120), .CO(n730), .S(n731) );
  CFA1X1 U574 ( .A(n1613), .B(n1090), .CI(n1036), .CO(n732), .S(n733) );
  CFA1X1 U575 ( .A(n952), .B(n1062), .CI(n1012), .CO(n734), .S(n735) );
  CHA1X1 U576 ( .A(n857), .B(n990), .CO(n736), .S(n737) );
  CFA1X1 U577 ( .A(n743), .B(n741), .CI(n754), .CO(n738), .S(n739) );
  CFA1X1 U578 ( .A(n758), .B(n756), .CI(n745), .CO(n740), .S(n741) );
  CFA1X1 U579 ( .A(n751), .B(n747), .CI(n749), .CO(n742), .S(n743) );
  CFA1X1 U580 ( .A(n764), .B(n762), .CI(n760), .CO(n744), .S(n745) );
  CFA1X1 U581 ( .A(n1013), .B(n1121), .CI(n1037), .CO(n746), .S(n747) );
  CFA1X1 U582 ( .A(n991), .B(n1091), .CI(n1063), .CO(n748), .S(n749) );
  CFA1X1 U583 ( .A(n1559), .B(n971), .CI(n953), .CO(n750), .S(n751) );
  CFA1X1 U584 ( .A(n757), .B(n755), .CI(n768), .CO(n752), .S(n753) );
  CFA1X1 U585 ( .A(n772), .B(n759), .CI(n770), .CO(n754), .S(n755) );
  CFA1X1 U586 ( .A(n774), .B(n761), .CI(n763), .CO(n756), .S(n757) );
  CFA1X1 U587 ( .A(n992), .B(n776), .CI(n765), .CO(n758), .S(n759) );
  CFA1X1 U588 ( .A(n954), .B(n1672), .CI(n1038), .CO(n760), .S(n761) );
  CFA1X1 U589 ( .A(n972), .B(n1561), .CI(n1122), .CO(n762), .S(n763) );
  CHA1X1 U590 ( .A(n858), .B(n1014), .CO(n764), .S(n765) );
  CFA1X1 U591 ( .A(n771), .B(n769), .CI(n780), .CO(n766), .S(n767) );
  CFA1X1 U592 ( .A(n775), .B(n782), .CI(n773), .CO(n768), .S(n769) );
  CFA1X1 U593 ( .A(n784), .B(n777), .CI(n786), .CO(n770), .S(n771) );
  CFA1X1 U594 ( .A(n1039), .B(n788), .CI(n1123), .CO(n772), .S(n773) );
  CFA1X1 U595 ( .A(n1015), .B(n1065), .CI(n1093), .CO(n774), .S(n775) );
  CFA1X1 U597 ( .A(n783), .B(n781), .CI(n792), .CO(n778), .S(n779) );
  CFA1X1 U598 ( .A(n787), .B(n794), .CI(n785), .CO(n780), .S(n781) );
  CFA1X1 U599 ( .A(n789), .B(n796), .CI(n798), .CO(n782), .S(n783) );
  CFA1X1 U600 ( .A(n994), .B(n1040), .CI(n1016), .CO(n784), .S(n785) );
  CFA1X1 U601 ( .A(n974), .B(n1066), .CI(n1124), .CO(n786), .S(n787) );
  CHA1X1 U602 ( .A(n859), .B(n1094), .CO(n788), .S(n789) );
  CFA1X1 U603 ( .A(n802), .B(n793), .CI(n795), .CO(n790), .S(n791) );
  CFA1X1 U604 ( .A(n799), .B(n804), .CI(n797), .CO(n792), .S(n793) );
  CFA1X1 U605 ( .A(n1125), .B(n806), .CI(n808), .CO(n794), .S(n795) );
  CFA1X1 U606 ( .A(n1095), .B(n1041), .CI(n1067), .CO(n796), .S(n797) );
  CFA1X1 U607 ( .A(n975), .B(n1017), .CI(n1623), .CO(n798), .S(n799) );
  CFA1X1 U608 ( .A(n805), .B(n803), .CI(n812), .CO(n800), .S(n801) );
  CFA1X1 U609 ( .A(n816), .B(n807), .CI(n814), .CO(n802), .S(n803) );
  CFA1X1 U610 ( .A(n1018), .B(n809), .CI(n1042), .CO(n804), .S(n805) );
  CFA1X1 U611 ( .A(n1625), .B(n1068), .CI(n1126), .CO(n806), .S(n807) );
  CHA1X1 U612 ( .A(n860), .B(n1096), .CO(n808), .S(n809) );
  CFA1X1 U613 ( .A(n815), .B(n813), .CI(n820), .CO(n810), .S(n811) );
  CFA1X1 U614 ( .A(n824), .B(n817), .CI(n822), .CO(n812), .S(n813) );
  CFA1X1 U615 ( .A(n1127), .B(n1097), .CI(n1069), .CO(n814), .S(n815) );
  CFA1X1 U617 ( .A(n828), .B(n821), .CI(n823), .CO(n818), .S(n819) );
  CFA1X1 U618 ( .A(n1044), .B(n830), .CI(n825), .CO(n820), .S(n821) );
  CFA1X1 U619 ( .A(n1020), .B(n1070), .CI(n1128), .CO(n822), .S(n823) );
  CHA1X1 U620 ( .A(n861), .B(n1098), .CO(n824), .S(n825) );
  CFA1X1 U621 ( .A(n834), .B(n829), .CI(n831), .CO(n826), .S(n827) );
  CFA1X1 U622 ( .A(n1099), .B(n836), .CI(n1071), .CO(n828), .S(n829) );
  CFA1X1 U623 ( .A(n1021), .B(n1129), .CI(n1045), .CO(n830), .S(n831) );
  CFA1X1 U624 ( .A(n837), .B(n835), .CI(n840), .CO(n832), .S(n833) );
  CFA1X1 U625 ( .A(n1630), .B(n1072), .CI(n1130), .CO(n834), .S(n835) );
  CHA1X1 U626 ( .A(n862), .B(n1100), .CO(n836), .S(n837) );
  CFA1X1 U627 ( .A(n1073), .B(n841), .CI(n844), .CO(n838), .S(n839) );
  CFA1X1 U629 ( .A(n1102), .B(n845), .CI(n1074), .CO(n842), .S(n843) );
  CHA1X1 U630 ( .A(n1132), .B(n863), .CO(n844), .S(n845) );
  CFA1X1 U631 ( .A(n1075), .B(n1103), .CI(n1133), .CO(n846), .S(n847) );
  CHA1X1 U632 ( .A(n1134), .B(n1104), .CO(n848), .S(n849) );
  COND2X1 U633 ( .A(n115), .B(n1468), .C(n114), .D(n1139), .Z(n850) );
  CND2IX1 U638 ( .B(n1736), .A(n113), .Z(n1139) );
  COND2X1 U639 ( .A(n112), .B(n1469), .C(n110), .D(n1144), .Z(n851) );
  COND2X1 U641 ( .A(n112), .B(n1142), .C(n110), .D(n1141), .Z(n869) );
  COND2X1 U653 ( .A(n107), .B(n1149), .C(n105), .D(n1148), .Z(n875) );
  COND2X1 U654 ( .A(n1150), .B(n107), .C(n105), .D(n1149), .Z(n876) );
  COND2X1 U663 ( .A(n102), .B(n1604), .C(n100), .D(n1160), .Z(n853) );
  COND2X1 U667 ( .A(n102), .B(n1156), .C(n100), .D(n1155), .Z(n881) );
  COND2X1 U681 ( .A(n97), .B(n1579), .C(n95), .D(n1171), .Z(n854) );
  COND2X1 U683 ( .A(n97), .B(n1163), .C(n1162), .D(n95), .Z(n887) );
  COND2X1 U686 ( .A(n97), .B(n1166), .C(n95), .D(n1165), .Z(n890) );
  COND2X1 U687 ( .A(n97), .B(n1167), .C(n95), .D(n1166), .Z(n891) );
  COND2X1 U688 ( .A(n97), .B(n1168), .C(n95), .D(n1167), .Z(n892) );
  COND2X1 U689 ( .A(n97), .B(n1169), .C(n95), .D(n1168), .Z(n893) );
  COND2X1 U703 ( .A(n91), .B(n1473), .C(n89), .D(n1184), .Z(n855) );
  COND2X1 U708 ( .A(n91), .B(n1177), .C(n1176), .D(n89), .Z(n900) );
  COND2X1 U709 ( .A(n91), .B(n1178), .C(n1177), .D(n89), .Z(n901) );
  COND2X1 U712 ( .A(n91), .B(n1181), .C(n1180), .D(n89), .Z(n904) );
  COND2X1 U714 ( .A(n1183), .B(n91), .C(n1182), .D(n89), .Z(n906) );
  COND2X1 U736 ( .A(n85), .B(n1192), .C(n1191), .D(n1566), .Z(n914) );
  COND2X1 U737 ( .A(n85), .B(n1193), .C(n1192), .D(n1627), .Z(n915) );
  COND2X1 U738 ( .A(n85), .B(n1194), .C(n1193), .D(n1566), .Z(n916) );
  COND2X1 U739 ( .A(n85), .B(n1195), .C(n1194), .D(n1566), .Z(n917) );
  COND2X1 U740 ( .A(n85), .B(n1196), .C(n1195), .D(n1566), .Z(n918) );
  COND2X1 U742 ( .A(n1198), .B(n85), .C(n1197), .D(n1566), .Z(n920) );
  CND2IX1 U758 ( .B(n1736), .A(n1697), .Z(n1199) );
  COND2X1 U766 ( .A(n77), .B(n1207), .C(n1206), .D(n74), .Z(n928) );
  COND2X1 U772 ( .A(n77), .B(n1213), .C(n1212), .D(n74), .Z(n934) );
  COND2X1 U798 ( .A(n69), .B(n1222), .C(n1221), .D(n66), .Z(n942) );
  COND2X1 U799 ( .A(n69), .B(n1223), .C(n1222), .D(n66), .Z(n943) );
  COND2X1 U801 ( .A(n69), .B(n1225), .C(n1224), .D(n66), .Z(n945) );
  COND2X1 U803 ( .A(n69), .B(n1227), .C(n1226), .D(n66), .Z(n947) );
  COND2X1 U804 ( .A(n69), .B(n1228), .C(n1227), .D(n66), .Z(n948) );
  COND2X1 U805 ( .A(n69), .B(n1229), .C(n1228), .D(n66), .Z(n949) );
  COND2X1 U809 ( .A(n69), .B(n1233), .C(n1232), .D(n66), .Z(n953) );
  COND2X1 U810 ( .A(n69), .B(n1234), .C(n1233), .D(n66), .Z(n954) );
  COND2X1 U838 ( .A(n61), .B(n1243), .C(n1242), .D(n58), .Z(n962) );
  COND2X1 U839 ( .A(n61), .B(n1244), .C(n1243), .D(n58), .Z(n963) );
  CND2IX1 U872 ( .B(n1736), .A(n1733), .Z(n1256) );
  COND2X1 U881 ( .A(n53), .B(n1265), .C(n1264), .D(n50), .Z(n983) );
  COND2X1 U884 ( .A(n53), .B(n1268), .C(n1267), .D(n50), .Z(n986) );
  COND2X1 U886 ( .A(n53), .B(n1270), .C(n1269), .D(n50), .Z(n988) );
  COND2X1 U889 ( .A(n53), .B(n1273), .C(n1272), .D(n50), .Z(n991) );
  CND2IX1 U918 ( .B(n1736), .A(n1730), .Z(n1279) );
  COND2X1 U923 ( .A(n44), .B(n1284), .C(n1283), .D(n42), .Z(n1001) );
  COND2X1 U925 ( .A(n44), .B(n1286), .C(n1285), .D(n42), .Z(n1003) );
  COND2X1 U926 ( .A(n44), .B(n1287), .C(n1286), .D(n42), .Z(n1004) );
  COND2X1 U928 ( .A(n44), .B(n1289), .C(n1288), .D(n42), .Z(n1006) );
  COND2X1 U929 ( .A(n44), .B(n1290), .C(n1289), .D(n42), .Z(n1007) );
  COND2X1 U931 ( .A(n44), .B(n1292), .C(n1291), .D(n42), .Z(n1009) );
  COND2X1 U932 ( .A(n44), .B(n1293), .C(n1292), .D(n42), .Z(n1010) );
  COND2X1 U934 ( .A(n44), .B(n1295), .C(n1294), .D(n42), .Z(n1012) );
  COND2X1 U935 ( .A(n44), .B(n1296), .C(n1295), .D(n42), .Z(n1013) );
  COND2X1 U936 ( .A(n44), .B(n1297), .C(n1296), .D(n42), .Z(n1014) );
  COND2X1 U937 ( .A(n44), .B(n1298), .C(n1297), .D(n42), .Z(n1015) );
  COND2X1 U938 ( .A(n44), .B(n1299), .C(n1298), .D(n42), .Z(n1016) );
  COND2X1 U939 ( .A(n44), .B(n1300), .C(n1299), .D(n42), .Z(n1017) );
  COND2X1 U941 ( .A(n44), .B(n1302), .C(n1301), .D(n42), .Z(n1019) );
  CND2IX1 U968 ( .B(n1736), .A(n1723), .Z(n1304) );
  COND2X1 U976 ( .A(n36), .B(n1312), .C(n1311), .D(n1679), .Z(n1028) );
  COND2X1 U977 ( .A(n36), .B(n1313), .C(n1312), .D(n1679), .Z(n1029) );
  COND2X1 U980 ( .A(n36), .B(n1316), .C(n1315), .D(n1679), .Z(n1032) );
  COND2X1 U982 ( .A(n36), .B(n1318), .C(n1317), .D(n1679), .Z(n1034) );
  COND2X1 U984 ( .A(n36), .B(n1320), .C(n1319), .D(n1679), .Z(n1036) );
  COND2X1 U985 ( .A(n36), .B(n1321), .C(n1320), .D(n1679), .Z(n1037) );
  COND2X1 U986 ( .A(n36), .B(n1322), .C(n1321), .D(n1679), .Z(n1038) );
  CND2IX1 U1022 ( .B(n1736), .A(n1718), .Z(n1331) );
  COND2X1 U1036 ( .A(n27), .B(n1345), .C(n1649), .D(n1344), .Z(n1060) );
  COND2X1 U1039 ( .A(n27), .B(n1348), .C(n1649), .D(n1347), .Z(n1063) );
  COND2X1 U1091 ( .A(n18), .B(n1371), .C(n1670), .D(n1370), .Z(n1085) );
  COND2X1 U1093 ( .A(n18), .B(n1373), .C(n1670), .D(n1372), .Z(n1087) );
  COND2X1 U1094 ( .A(n18), .B(n1374), .C(n1670), .D(n1373), .Z(n1088) );
  COND2X1 U1097 ( .A(n18), .B(n1377), .C(n1670), .D(n1376), .Z(n1091) );
  CND2IX1 U1142 ( .B(n1736), .A(n1637), .Z(n1391) );
  COND2X1 U1144 ( .A(n9), .B(n1393), .C(n1564), .D(n1392), .Z(n1106) );
  COND2X1 U1145 ( .A(n9), .B(n1394), .C(n1564), .D(n1393), .Z(n1107) );
  COND2X1 U1146 ( .A(n9), .B(n1395), .C(n1564), .D(n1394), .Z(n1108) );
  COND2X1 U1147 ( .A(n9), .B(n1396), .C(n1564), .D(n1395), .Z(n1109) );
  COND2X1 U1149 ( .A(n9), .B(n1398), .C(n1564), .D(n1397), .Z(n1111) );
  COND2X1 U1150 ( .A(n9), .B(n1399), .C(n1564), .D(n1398), .Z(n1112) );
  COND2X1 U1152 ( .A(n9), .B(n1401), .C(n1564), .D(n1400), .Z(n1114) );
  COND2X1 U1153 ( .A(n9), .B(n1402), .C(n1564), .D(n1401), .Z(n1115) );
  COND2X1 U1154 ( .A(n9), .B(n1403), .C(n1564), .D(n1402), .Z(n1116) );
  COND2X1 U1155 ( .A(n9), .B(n1404), .C(n1564), .D(n1403), .Z(n1117) );
  COND2X1 U1157 ( .A(n9), .B(n1406), .C(n1564), .D(n1405), .Z(n1119) );
  COND2X1 U1158 ( .A(n9), .B(n1407), .C(n1564), .D(n1406), .Z(n1120) );
  COND2X1 U1159 ( .A(n9), .B(n1408), .C(n1564), .D(n1407), .Z(n1121) );
  COND2X1 U1160 ( .A(n9), .B(n1409), .C(n1564), .D(n1408), .Z(n1122) );
  COND2X1 U1161 ( .A(n9), .B(n1410), .C(n1564), .D(n1409), .Z(n1123) );
  COND2X1 U1163 ( .A(n9), .B(n1412), .C(n1564), .D(n1411), .Z(n1125) );
  COND2X1 U1164 ( .A(n9), .B(n1413), .C(n1564), .D(n1412), .Z(n1126) );
  COND2X1 U1165 ( .A(n9), .B(n1414), .C(n1564), .D(n1413), .Z(n1127) );
  COND2X1 U1166 ( .A(n9), .B(n1415), .C(n1564), .D(n1414), .Z(n1128) );
  COND2X1 U1167 ( .A(n9), .B(n1416), .C(n1564), .D(n1415), .Z(n1129) );
  COND2X1 U1168 ( .A(n9), .B(n1417), .C(n1564), .D(n1416), .Z(n1130) );
  COND2X1 U1169 ( .A(n9), .B(n1418), .C(n1564), .D(n1417), .Z(n1131) );
  COND2X1 U1170 ( .A(n9), .B(n1419), .C(n1564), .D(n1418), .Z(n1132) );
  COND2X1 U1171 ( .A(n9), .B(n1420), .C(n1564), .D(n1419), .Z(n1133) );
  COND2X1 U1172 ( .A(n9), .B(n1421), .C(n1564), .D(n1420), .Z(n1134) );
  COND2X1 U1173 ( .A(n9), .B(n1422), .C(n1564), .D(n1421), .Z(n1135) );
  COND2X1 U1174 ( .A(n9), .B(n1423), .C(n1564), .D(n1422), .Z(n1136) );
  CND2IX1 U1208 ( .B(n1736), .A(n1631), .Z(n1424) );
  CIVDX1 U1281 ( .A(n82), .Z0(n1565), .Z1(n1566) );
  CENX2 U1282 ( .A(n1696), .B(a[18]), .Z(n82) );
  COND2X1 U1283 ( .A(n85), .B(n1190), .C(n1189), .D(n1566), .Z(n912) );
  CNR2X1 U1284 ( .A(n53), .B(n1262), .Z(n1645) );
  CENX1 U1285 ( .A(n1697), .B(n1681), .Z(n1196) );
  CENXL U1286 ( .A(n1696), .B(n1681), .Z(n1213) );
  CENXL U1287 ( .A(n1695), .B(n1681), .Z(n1232) );
  CNIVX3 U1288 ( .A(n87), .Z(n1698) );
  CND2X2 U1289 ( .A(n1446), .B(n100), .Z(n102) );
  CND3X2 U1290 ( .A(n1598), .B(n1599), .C(n1600), .Z(n544) );
  CIVXL U1291 ( .A(n217), .Z(n1557) );
  CIVXL U1292 ( .A(n1557), .Z(n1558) );
  COND2X1 U1293 ( .A(n69), .B(n1226), .C(n1225), .D(n66), .Z(n946) );
  CENXL U1294 ( .A(n1695), .B(n1688), .Z(n1225) );
  CNIVX8 U1295 ( .A(n120), .Z(n1680) );
  CENXL U1296 ( .A(n1714), .B(n1682), .Z(n1356) );
  CENXL U1297 ( .A(n1631), .B(n1682), .Z(n1420) );
  CENXL U1298 ( .A(n1724), .B(n1682), .Z(n1300) );
  CENXL U1299 ( .A(n1695), .B(n1682), .Z(n1231) );
  CENXL U1300 ( .A(n1682), .B(n1700), .Z(n1156) );
  CENX1 U1301 ( .A(n1732), .B(n1682), .Z(n1252) );
  CND2X1 U1302 ( .A(n1700), .B(a[26]), .Z(n1606) );
  CND2X4 U1303 ( .A(n1639), .B(n1640), .Z(n1649) );
  CNIVX8 U1304 ( .A(n128), .Z(n1684) );
  CEOX2 U1305 ( .A(a[4]), .B(n1713), .Z(n1456) );
  CNIVX2 U1306 ( .A(n93), .Z(n1699) );
  CND2X2 U1307 ( .A(n391), .B(n1655), .Z(n245) );
  CNIVX1 U1308 ( .A(n937), .Z(n1559) );
  CIVX4 U1309 ( .A(n1633), .Z(n1634) );
  CENXL U1310 ( .A(n1695), .B(n1686), .Z(n1227) );
  COND2X1 U1311 ( .A(n61), .B(n1254), .C(n1253), .D(n58), .Z(n973) );
  CENX1 U1312 ( .A(n1732), .B(n1681), .Z(n1253) );
  CFA1X2 U1313 ( .A(n928), .B(n1082), .CI(n944), .CO(n580), .S(n581) );
  CFA1XL U1314 ( .A(n911), .B(n1025), .CI(n925), .CO(n506), .S(n507) );
  COND2XL U1315 ( .A(n44), .B(n1281), .C(n1280), .D(n42), .Z(n998) );
  COND2XL U1316 ( .A(n44), .B(n1294), .C(n1293), .D(n42), .Z(n1011) );
  COND2XL U1317 ( .A(n44), .B(n1291), .C(n1290), .D(n42), .Z(n1008) );
  COND2XL U1318 ( .A(n44), .B(n1288), .C(n1287), .D(n42), .Z(n1005) );
  COND2XL U1319 ( .A(n44), .B(n1301), .C(n1300), .D(n42), .Z(n1018) );
  COND2XL U1320 ( .A(n44), .B(n1582), .C(n1304), .D(n42), .Z(n861) );
  COND2XL U1321 ( .A(n44), .B(n1285), .C(n1284), .D(n42), .Z(n1002) );
  COND2X1 U1322 ( .A(n27), .B(n1337), .C(n1649), .D(n1336), .Z(n1052) );
  CENXL U1323 ( .A(n1712), .B(n156), .Z(n1337) );
  CENXL U1324 ( .A(n1732), .B(n1689), .Z(n1245) );
  CENXL U1325 ( .A(n1732), .B(n1688), .Z(n1246) );
  CENXL U1326 ( .A(n1732), .B(n1684), .Z(n1250) );
  CENXL U1327 ( .A(n1732), .B(n1691), .Z(n1243) );
  CENXL U1328 ( .A(n1732), .B(n1690), .Z(n1244) );
  CENXL U1329 ( .A(n1732), .B(n1685), .Z(n1249) );
  CENXL U1330 ( .A(n1732), .B(n1680), .Z(n1254) );
  CND2X2 U1331 ( .A(n1451), .B(n66), .Z(n69) );
  CIVXL U1332 ( .A(n1064), .Z(n1560) );
  CIVX2 U1333 ( .A(n1560), .Z(n1561) );
  CENXL U1334 ( .A(n1712), .B(n155), .Z(n1338) );
  CENX1 U1335 ( .A(n1631), .B(n152), .Z(n1405) );
  CENX1 U1336 ( .A(n1725), .B(n152), .Z(n1285) );
  CENXL U1337 ( .A(n1721), .B(n152), .Z(n1312) );
  COND2X1 U1338 ( .A(n77), .B(n1208), .C(n1207), .D(n74), .Z(n929) );
  CENXL U1339 ( .A(n1696), .B(n1686), .Z(n1208) );
  CFA1X2 U1340 ( .A(n1004), .B(n1112), .CI(n1028), .CO(n576), .S(n577) );
  CIVXL U1341 ( .A(a[10]), .Z(n1583) );
  CENXL U1342 ( .A(a[10]), .B(n1730), .Z(n1650) );
  COND2XL U1343 ( .A(n27), .B(n1357), .C(n1649), .D(n1356), .Z(n1072) );
  COND2XL U1344 ( .A(n27), .B(n1347), .C(n1649), .D(n1346), .Z(n1062) );
  COND2XL U1345 ( .A(n27), .B(n1352), .C(n1649), .D(n1351), .Z(n1067) );
  COND2XL U1346 ( .A(n27), .B(n1339), .C(n1649), .D(n1338), .Z(n1054) );
  COND2XL U1347 ( .A(n27), .B(n1349), .C(n1649), .D(n1348), .Z(n1064) );
  CND2X4 U1348 ( .A(n1456), .B(n1649), .Z(n27) );
  CIVXL U1349 ( .A(n352), .Z(n351) );
  COND1X1 U1350 ( .A(n352), .B(n340), .C(n341), .Z(n339) );
  CIVX2 U1351 ( .A(n1669), .Z(n1670) );
  CEOX2 U1352 ( .A(n1703), .B(a[2]), .Z(n1669) );
  CENXL U1353 ( .A(n1698), .B(n1690), .Z(n1172) );
  CENXL U1354 ( .A(n1681), .B(n1698), .Z(n1181) );
  CENXL U1355 ( .A(n1735), .B(n1698), .Z(n1183) );
  CENXL U1356 ( .A(n1698), .B(n1688), .Z(n1174) );
  CENXL U1357 ( .A(n1698), .B(n1689), .Z(n1173) );
  CENXL U1358 ( .A(n1698), .B(n1687), .Z(n1175) );
  CENXL U1359 ( .A(n1698), .B(n1686), .Z(n1176) );
  CENXL U1360 ( .A(n1682), .B(n1698), .Z(n1180) );
  CENXL U1361 ( .A(n1698), .B(n1685), .Z(n1177) );
  CENXL U1362 ( .A(n1680), .B(n1698), .Z(n1182) );
  CENXL U1363 ( .A(n1684), .B(n1698), .Z(n1178) );
  CENXL U1364 ( .A(n1683), .B(n1698), .Z(n1179) );
  CEOX1 U1365 ( .A(a[20]), .B(n1698), .Z(n1448) );
  CIVX3 U1366 ( .A(n1734), .Z(n1732) );
  CND2X2 U1367 ( .A(n1454), .B(n42), .Z(n44) );
  CEOX1 U1368 ( .A(a[8]), .B(n1727), .Z(n1454) );
  CIVX4 U1369 ( .A(n1668), .Z(n42) );
  COR2XL U1370 ( .A(n1196), .B(n1627), .Z(n1636) );
  COR2XL U1371 ( .A(n85), .B(n1197), .Z(n1635) );
  CNIVX2 U1372 ( .A(n138), .Z(n1689) );
  CNIVX2 U1373 ( .A(n146), .Z(n1693) );
  CNIVX3 U1374 ( .A(n130), .Z(n1685) );
  CENX1 U1375 ( .A(n1712), .B(n154), .Z(n1339) );
  CNIVX2 U1376 ( .A(n132), .Z(n1686) );
  CNIVX2 U1377 ( .A(n148), .Z(n1694) );
  CEOX1 U1378 ( .A(n1634), .B(n1695), .Z(n1451) );
  CANR1XL U1379 ( .A(n348), .B(n1661), .C(n343), .Z(n341) );
  CENX1 U1380 ( .A(n1735), .B(n1714), .Z(n1359) );
  CND2X1 U1381 ( .A(n587), .B(n608), .Z(n250) );
  CND2X1 U1382 ( .A(n631), .B(n650), .Z(n270) );
  CENX1 U1383 ( .A(n1695), .B(n1683), .Z(n1230) );
  CENX1 U1384 ( .A(n1695), .B(n1684), .Z(n1229) );
  CENX1 U1385 ( .A(n1708), .B(n152), .Z(n1372) );
  CENX1 U1386 ( .A(n1695), .B(n1685), .Z(n1228) );
  CENX1 U1387 ( .A(n1696), .B(n1684), .Z(n1210) );
  CENX1 U1388 ( .A(n1696), .B(n1685), .Z(n1209) );
  CENX1 U1389 ( .A(n1697), .B(n1683), .Z(n1194) );
  CENX1 U1390 ( .A(n1735), .B(n1699), .Z(n1170) );
  CENX1 U1391 ( .A(n1695), .B(n1680), .Z(n1233) );
  CENX1 U1392 ( .A(n1736), .B(n1695), .Z(n1234) );
  CENX1 U1393 ( .A(n1736), .B(n1696), .Z(n1215) );
  CENX1 U1394 ( .A(n1718), .B(n1692), .Z(n1317) );
  CND2X1 U1395 ( .A(n1635), .B(n1636), .Z(n919) );
  CENX1 U1396 ( .A(n1681), .B(n1700), .Z(n1157) );
  CENX1 U1397 ( .A(n1683), .B(n1699), .Z(n1166) );
  CENX1 U1398 ( .A(n1695), .B(n1691), .Z(n1222) );
  CENX1 U1399 ( .A(n1682), .B(n1699), .Z(n1167) );
  CENX1 U1400 ( .A(n1681), .B(n1699), .Z(n1168) );
  CENX1 U1401 ( .A(n1680), .B(n1699), .Z(n1169) );
  CENX1 U1402 ( .A(n1695), .B(n1687), .Z(n1226) );
  CENX1 U1403 ( .A(n1684), .B(n1699), .Z(n1165) );
  CENX1 U1404 ( .A(n1697), .B(n1689), .Z(n1188) );
  CNIVX2 U1405 ( .A(n142), .Z(n1691) );
  CIVX2 U1406 ( .A(n55), .Z(n1734) );
  CENX1 U1407 ( .A(n1685), .B(n1699), .Z(n1164) );
  CENX1 U1408 ( .A(n1696), .B(n1691), .Z(n1203) );
  CENX1 U1409 ( .A(n1730), .B(n152), .Z(n1260) );
  CENX1 U1410 ( .A(n1695), .B(n1693), .Z(n1220) );
  CNIVX1 U1411 ( .A(n960), .Z(n1619) );
  CENX1 U1412 ( .A(n1705), .B(n157), .Z(n1367) );
  CENX1 U1413 ( .A(n1695), .B(n1689), .Z(n1224) );
  CENX1 U1414 ( .A(n1695), .B(n1690), .Z(n1223) );
  CENX1 U1415 ( .A(n1696), .B(n1687), .Z(n1207) );
  CNIVX1 U1416 ( .A(n884), .Z(n1618) );
  CENX1 U1417 ( .A(n1735), .B(n1727), .Z(n1303) );
  CNIVX2 U1418 ( .A(n136), .Z(n1688) );
  CENX1 U1419 ( .A(n1684), .B(n1700), .Z(n1154) );
  CENX1 U1420 ( .A(n1686), .B(n1699), .Z(n1163) );
  CND2IX2 U1421 ( .B(n1650), .A(n50), .Z(n53) );
  CIVX3 U1422 ( .A(n1734), .Z(n1733) );
  CENX1 U1423 ( .A(n1695), .B(n1694), .Z(n1219) );
  CENX1 U1424 ( .A(n1733), .B(n152), .Z(n1237) );
  CNIVX3 U1425 ( .A(n126), .Z(n1683) );
  CNIVX2 U1426 ( .A(n124), .Z(n1682) );
  CNIVX2 U1427 ( .A(n122), .Z(n1681) );
  CEOX1 U1428 ( .A(a[6]), .B(n1721), .Z(n1455) );
  CNIVX2 U1429 ( .A(n33), .Z(n1679) );
  CENX1 U1430 ( .A(n1724), .B(n157), .Z(n1280) );
  CENX1 U1431 ( .A(n1688), .B(n1699), .Z(n1161) );
  CND2X2 U1432 ( .A(n95), .B(n1447), .Z(n97) );
  CND2X1 U1433 ( .A(n1580), .B(n1581), .Z(n1447) );
  CENX2 U1434 ( .A(n1698), .B(a[22]), .Z(n95) );
  CENX1 U1435 ( .A(n1687), .B(n1699), .Z(n1162) );
  CENX1 U1436 ( .A(n1686), .B(n1700), .Z(n1152) );
  CENX1 U1437 ( .A(n1695), .B(n151), .Z(n1217) );
  CENX1 U1438 ( .A(n1696), .B(n1694), .Z(n1200) );
  CND2X1 U1439 ( .A(n1711), .B(n1638), .Z(n1640) );
  CNIVX1 U1440 ( .A(n116), .Z(n1735) );
  CANR1XL U1441 ( .A(n1662), .B(n357), .C(n354), .Z(n352) );
  CANR1X1 U1442 ( .A(n288), .B(n1657), .C(n283), .Z(n281) );
  CANR1XL U1443 ( .A(n381), .B(n1665), .C(n378), .Z(n376) );
  COND1XL U1444 ( .A(n328), .B(n322), .C(n323), .Z(n321) );
  CNIVX1 U1445 ( .A(n116), .Z(n1736) );
  CND2X1 U1446 ( .A(n539), .B(n562), .Z(n235) );
  CANR1XL U1447 ( .A(n365), .B(n1666), .C(n362), .Z(n360) );
  CENX1 U1448 ( .A(n251), .B(n173), .Z(product[24]) );
  CENX1 U1449 ( .A(n271), .B(n175), .Z(product[22]) );
  CENX1 U1450 ( .A(n304), .B(n180), .Z(product[17]) );
  CENX1 U1451 ( .A(n297), .B(n179), .Z(product[18]) );
  CENX1 U1452 ( .A(n191), .B(n365), .Z(product[6]) );
  CENX1 U1453 ( .A(n260), .B(n174), .Z(product[23]) );
  CENXL U1454 ( .A(n1716), .B(n1694), .Z(n1344) );
  CNIVX3 U1455 ( .A(n99), .Z(n1700) );
  CNIVX3 U1456 ( .A(n1702), .Z(n1631) );
  CIVX2 U1457 ( .A(n1711), .Z(n1707) );
  CIVX1 U1458 ( .A(n1717), .Z(n1714) );
  CIVX2 U1459 ( .A(n1722), .Z(n1721) );
  COAN1XL U1460 ( .A(n330), .B(n313), .C(n314), .Z(n1562) );
  CIVX2 U1461 ( .A(n1700), .Z(n1604) );
  CIVDX3 U1462 ( .A(n1628), .Z0(n1563), .Z1(n1564) );
  CNIVX1 U1463 ( .A(n12), .Z(n1637) );
  CIVX2 U1464 ( .A(n1704), .Z(n1702) );
  COR2X1 U1465 ( .A(n631), .B(n650), .Z(n1567) );
  COND2X1 U1466 ( .A(n85), .B(n1191), .C(n1190), .D(n1627), .Z(n913) );
  COND2X1 U1467 ( .A(n107), .B(n1147), .C(n105), .D(n1146), .Z(n873) );
  COR2XL U1468 ( .A(n539), .B(n562), .Z(n1568) );
  CIVX2 U1469 ( .A(n1699), .Z(n1579) );
  CNIVX4 U1470 ( .A(n63), .Z(n1695) );
  CIVX2 U1471 ( .A(n1695), .Z(n1586) );
  COR2X1 U1472 ( .A(n1136), .B(n865), .Z(n1569) );
  CND2X4 U1473 ( .A(n89), .B(n1448), .Z(n91) );
  COND2X1 U1474 ( .A(n1151), .B(n105), .C(n1470), .D(n107), .Z(n852) );
  CENX1 U1475 ( .A(n1683), .B(n1700), .Z(n1155) );
  CFA1XL U1476 ( .A(n946), .B(n1056), .CI(n1006), .CO(n622), .S(n623) );
  CENXL U1477 ( .A(n1729), .B(n154), .Z(n1258) );
  CENXL U1478 ( .A(n1695), .B(n150), .Z(n1218) );
  CENXL U1479 ( .A(n1695), .B(n1692), .Z(n1221) );
  CENX1 U1480 ( .A(n1696), .B(n1688), .Z(n1206) );
  CENX1 U1481 ( .A(n1696), .B(n1689), .Z(n1205) );
  COND2X1 U1482 ( .A(n27), .B(n1346), .C(n1649), .D(n1345), .Z(n1061) );
  COND2X1 U1483 ( .A(n27), .B(n1338), .C(n1649), .D(n1337), .Z(n1053) );
  CNIVX1 U1484 ( .A(n930), .Z(n1570) );
  CFA1X1 U1485 ( .A(n904), .B(n984), .CI(n1570), .CO(n626), .S(n627) );
  CNR2IX1 U1486 ( .B(n1736), .A(n110), .Z(n871) );
  COND2XL U1487 ( .A(n1143), .B(n112), .C(n110), .D(n1142), .Z(n870) );
  COND2XL U1488 ( .A(n112), .B(n1141), .C(n110), .D(n1140), .Z(n868) );
  CENX1 U1489 ( .A(n1701), .B(a[28]), .Z(n110) );
  CND2XL U1490 ( .A(n385), .B(n207), .Z(n167) );
  CENX1 U1491 ( .A(n1706), .B(n155), .Z(n1369) );
  CND2IXL U1492 ( .B(n1736), .A(n1699), .Z(n1171) );
  CND2X1 U1493 ( .A(n1578), .B(n1699), .Z(n1581) );
  CFA1XL U1494 ( .A(n969), .B(n1061), .CI(n1119), .CO(n718), .S(n719) );
  COND2X1 U1495 ( .A(n61), .B(n1247), .C(n1246), .D(n58), .Z(n966) );
  CNR2XL U1496 ( .A(n539), .B(n562), .Z(n1571) );
  CND2IXL U1497 ( .B(n1736), .A(n1700), .Z(n1160) );
  CENXL U1498 ( .A(n1735), .B(n1700), .Z(n1159) );
  CENXL U1499 ( .A(n1685), .B(n1700), .Z(n1153) );
  CENXL U1500 ( .A(n1680), .B(n1700), .Z(n1158) );
  CEOX4 U1501 ( .A(n1563), .B(n1702), .Z(n1458) );
  COND2X1 U1502 ( .A(n91), .B(n1179), .C(n1178), .D(n89), .Z(n902) );
  COND2X1 U1503 ( .A(n9), .B(n1400), .C(n1564), .D(n1399), .Z(n1113) );
  COND2X1 U1504 ( .A(n1170), .B(n97), .C(n95), .D(n1169), .Z(n894) );
  CENX1 U1505 ( .A(n1632), .B(n153), .Z(n1404) );
  COND2X1 U1506 ( .A(n97), .B(n1165), .C(n1164), .D(n95), .Z(n889) );
  CFA1XL U1507 ( .A(n889), .B(n941), .CI(n899), .CO(n508), .S(n509) );
  COND2XL U1508 ( .A(n97), .B(n1164), .C(n1163), .D(n95), .Z(n888) );
  COND2X1 U1509 ( .A(n102), .B(n1158), .C(n100), .D(n1157), .Z(n883) );
  COND2X1 U1510 ( .A(n102), .B(n1155), .C(n100), .D(n1154), .Z(n880) );
  COND1X1 U1511 ( .A(n280), .B(n292), .C(n281), .Z(n1572) );
  COND1XL U1512 ( .A(n280), .B(n292), .C(n281), .Z(n279) );
  CIVXL U1513 ( .A(n239), .Z(n390) );
  CANR1X1 U1514 ( .A(n229), .B(n216), .C(n217), .Z(n1573) );
  CANR1XL U1515 ( .A(n229), .B(n216), .C(n1558), .Z(n215) );
  CHA1XL U1516 ( .A(n882), .B(n852), .CO(n536), .S(n537) );
  CEO3X2 U1517 ( .A(n582), .B(n576), .C(n580), .Z(n1574) );
  CENXL U1518 ( .A(n199), .B(n1575), .Z(product[31]) );
  CAN2X1 U1519 ( .A(n1663), .B(n198), .Z(n1575) );
  CENX1 U1520 ( .A(a[2]), .B(n1710), .Z(n1648) );
  COAN1X1 U1521 ( .A(n259), .B(n249), .C(n250), .Z(n246) );
  CIVDXL U1522 ( .A(n259), .Z0(n257) );
  CANR1X1 U1523 ( .A(n228), .B(n241), .C(n229), .Z(n227) );
  CENX4 U1524 ( .A(n1699), .B(a[24]), .Z(n100) );
  CND2X1 U1525 ( .A(n551), .B(n572), .Z(n1600) );
  CND2X1 U1526 ( .A(n574), .B(n551), .Z(n1598) );
  CANR1X2 U1527 ( .A(n243), .B(n1572), .C(n244), .Z(n1576) );
  COND1X2 U1528 ( .A(n262), .B(n245), .C(n246), .Z(n244) );
  CANR1X1 U1529 ( .A(n243), .B(n279), .C(n244), .Z(n242) );
  COND2X1 U1530 ( .A(n18), .B(n1381), .C(n1670), .D(n1380), .Z(n1095) );
  CIVX1 U1531 ( .A(n1092), .Z(n1671) );
  COND2X1 U1532 ( .A(n18), .B(n1378), .C(n1670), .D(n1377), .Z(n1092) );
  CND2X2 U1533 ( .A(n1445), .B(n105), .Z(n107) );
  CFA1X1 U1534 ( .A(n966), .B(n1086), .CI(n1116), .CO(n662), .S(n663) );
  COND2X1 U1535 ( .A(n18), .B(n1375), .C(n1670), .D(n1374), .Z(n1089) );
  CIVXL U1536 ( .A(n261), .Z(n263) );
  CND2X1 U1537 ( .A(n1567), .B(n394), .Z(n261) );
  CIVXL U1538 ( .A(n292), .Z(n291) );
  CIVXL U1539 ( .A(n322), .Z(n401) );
  COND2XL U1540 ( .A(n9), .B(n1405), .C(n1564), .D(n1404), .Z(n1118) );
  CFA1XL U1541 ( .A(n880), .B(n910), .CI(n851), .CO(n482), .S(n483) );
  COND1X1 U1542 ( .A(n358), .B(n360), .C(n359), .Z(n357) );
  COND2X1 U1543 ( .A(n27), .B(n1343), .C(n1649), .D(n1342), .Z(n1058) );
  CENXL U1544 ( .A(n1684), .B(n1701), .Z(n1145) );
  CND2IXL U1545 ( .B(n1736), .A(n1701), .Z(n1151) );
  CENXL U1546 ( .A(n1735), .B(n1701), .Z(n1150) );
  CENXL U1547 ( .A(n1682), .B(n1701), .Z(n1147) );
  CENXL U1548 ( .A(n1683), .B(n1701), .Z(n1146) );
  CENXL U1549 ( .A(n1680), .B(n1701), .Z(n1149) );
  CENXL U1550 ( .A(n1681), .B(n1701), .Z(n1148) );
  CEOX1 U1551 ( .A(a[26]), .B(n1701), .Z(n1445) );
  CNIVX4 U1552 ( .A(n71), .Z(n1696) );
  CFA1X1 U1553 ( .A(n906), .B(n1058), .CI(n986), .CO(n664), .S(n665) );
  CIVXL U1554 ( .A(n272), .Z(n394) );
  COND2X1 U1555 ( .A(n69), .B(n1231), .C(n1230), .D(n66), .Z(n951) );
  CFA1XL U1556 ( .A(n929), .B(n1083), .CI(n963), .CO(n602), .S(n603) );
  COND2X1 U1557 ( .A(n9), .B(n1411), .C(n1564), .D(n1410), .Z(n1124) );
  CFA1X1 U1558 ( .A(n967), .B(n1087), .CI(n1117), .CO(n682), .S(n683) );
  COND2X1 U1559 ( .A(n18), .B(n1372), .C(n1670), .D(n1371), .Z(n1086) );
  CNR2IX1 U1560 ( .B(n1736), .A(n1566), .Z(n921) );
  COND2X1 U1561 ( .A(n85), .B(n1189), .C(n1188), .D(n1566), .Z(n911) );
  CENXL U1562 ( .A(n167), .B(n1647), .Z(product[30]) );
  COND1XL U1563 ( .A(n214), .B(n1576), .C(n215), .Z(n1577) );
  COND1X1 U1564 ( .A(n214), .B(n242), .C(n1573), .Z(n213) );
  CIVXL U1565 ( .A(n229), .Z(n231) );
  COND1XL U1566 ( .A(n330), .B(n313), .C(n314), .Z(n312) );
  CIVXL U1567 ( .A(n330), .Z(n329) );
  CFA1XL U1568 ( .A(n897), .B(n977), .CI(n923), .CO(n452), .S(n453) );
  CIVX1 U1569 ( .A(n206), .Z(n385) );
  CNR2X2 U1570 ( .A(n431), .B(n458), .Z(n206) );
  CNR2X2 U1571 ( .A(n707), .B(n722), .Z(n295) );
  COND2X1 U1572 ( .A(n69), .B(n1232), .C(n1231), .D(n66), .Z(n952) );
  CND2X1 U1573 ( .A(a[22]), .B(n1579), .Z(n1580) );
  CIVXL U1574 ( .A(a[22]), .Z(n1578) );
  CND2XL U1575 ( .A(n39), .B(a[10]), .Z(n1584) );
  CND2X1 U1576 ( .A(n1582), .B(n1583), .Z(n1585) );
  CND2X2 U1577 ( .A(n1584), .B(n1585), .Z(n50) );
  CIVX2 U1578 ( .A(n39), .Z(n1582) );
  COND2XL U1579 ( .A(n53), .B(n1266), .C(n1265), .D(n50), .Z(n984) );
  COND2XL U1580 ( .A(n53), .B(n1267), .C(n1266), .D(n50), .Z(n985) );
  COND2X1 U1581 ( .A(n53), .B(n1259), .C(n1258), .D(n50), .Z(n977) );
  COND2X1 U1582 ( .A(n53), .B(n1275), .C(n1274), .D(n50), .Z(n993) );
  COND2X1 U1583 ( .A(n53), .B(n1263), .C(n1262), .D(n50), .Z(n981) );
  COND2X1 U1584 ( .A(n53), .B(n1272), .C(n1271), .D(n50), .Z(n990) );
  CND2XL U1585 ( .A(n1695), .B(a[16]), .Z(n1588) );
  CND2X1 U1586 ( .A(n1586), .B(n1587), .Z(n1589) );
  CND2X2 U1587 ( .A(n1588), .B(n1589), .Z(n74) );
  CIVX1 U1588 ( .A(a[16]), .Z(n1587) );
  COND2XL U1589 ( .A(n77), .B(n1212), .C(n1211), .D(n74), .Z(n933) );
  COND2XL U1590 ( .A(n77), .B(n1211), .C(n1210), .D(n74), .Z(n932) );
  COND2XL U1591 ( .A(n77), .B(n1210), .C(n1209), .D(n74), .Z(n931) );
  COND2XL U1592 ( .A(n77), .B(n1209), .C(n1208), .D(n74), .Z(n930) );
  COND2X1 U1593 ( .A(n77), .B(n1205), .C(n1204), .D(n74), .Z(n926) );
  COND2X1 U1594 ( .A(n77), .B(n1206), .C(n1205), .D(n74), .Z(n927) );
  COND2X1 U1595 ( .A(n77), .B(n1475), .C(n74), .D(n1216), .Z(n857) );
  CNR2IXL U1596 ( .B(n1736), .A(n74), .Z(n937) );
  CND2IX4 U1597 ( .B(n1651), .A(n74), .Z(n77) );
  CEOX2 U1598 ( .A(n635), .B(n652), .Z(n1590) );
  CEOX2 U1599 ( .A(n1590), .B(n633), .Z(n631) );
  CND2XL U1600 ( .A(n633), .B(n652), .Z(n1591) );
  CND2X1 U1601 ( .A(n633), .B(n635), .Z(n1592) );
  CND2XL U1602 ( .A(n652), .B(n635), .Z(n1593) );
  CND3X1 U1603 ( .A(n1591), .B(n1592), .C(n1593), .Z(n630) );
  CEO3X1 U1604 ( .A(n602), .B(n583), .C(n600), .Z(n573) );
  CND2X1 U1605 ( .A(n602), .B(n583), .Z(n1594) );
  CND2X1 U1606 ( .A(n602), .B(n600), .Z(n1595) );
  CND2X1 U1607 ( .A(n583), .B(n600), .Z(n1596) );
  CND3X2 U1608 ( .A(n1594), .B(n1595), .C(n1596), .Z(n572) );
  CEOX2 U1609 ( .A(n574), .B(n1574), .Z(n1597) );
  CEOX2 U1610 ( .A(n1597), .B(n572), .Z(n545) );
  CND2X1 U1611 ( .A(n574), .B(n572), .Z(n1599) );
  CND2X1 U1612 ( .A(a[24]), .B(n1604), .Z(n1602) );
  CND2XL U1613 ( .A(n1601), .B(n1700), .Z(n1603) );
  CND2X1 U1614 ( .A(n1602), .B(n1603), .Z(n1446) );
  CIVXL U1615 ( .A(a[24]), .Z(n1601) );
  CND2X1 U1616 ( .A(n1604), .B(n1605), .Z(n1607) );
  CND2X2 U1617 ( .A(n1606), .B(n1607), .Z(n105) );
  CIVX2 U1618 ( .A(a[26]), .Z(n1605) );
  COND2XL U1619 ( .A(n107), .B(n1146), .C(n105), .D(n1145), .Z(n872) );
  COND2XL U1620 ( .A(n107), .B(n1148), .C(n105), .D(n1147), .Z(n874) );
  CNR2IX1 U1621 ( .B(n1736), .A(n105), .Z(n877) );
  CEOX2 U1622 ( .A(n591), .B(n610), .Z(n1608) );
  CEOX2 U1623 ( .A(n1608), .B(n589), .Z(n587) );
  CND2XL U1624 ( .A(n589), .B(n610), .Z(n1609) );
  CND2X1 U1625 ( .A(n589), .B(n591), .Z(n1610) );
  CND2XL U1626 ( .A(n610), .B(n591), .Z(n1611) );
  CND3XL U1627 ( .A(n1609), .B(n1610), .C(n1611), .Z(n586) );
  CNIVX4 U1628 ( .A(n79), .Z(n1697) );
  CANR1XL U1629 ( .A(n1653), .B(n213), .C(n1676), .Z(n199) );
  CIVX2 U1630 ( .A(n1576), .Z(n241) );
  CENXL U1631 ( .A(n1577), .B(n168), .Z(product[29]) );
  CIVX1 U1632 ( .A(n936), .Z(n1612) );
  CIVX2 U1633 ( .A(n1612), .Z(n1613) );
  CIVXL U1634 ( .A(n1059), .Z(n1614) );
  CIVX1 U1635 ( .A(n1614), .Z(n1615) );
  CIVXL U1636 ( .A(n1057), .Z(n1616) );
  CIVX1 U1637 ( .A(n1616), .Z(n1617) );
  CENXL U1638 ( .A(n1682), .B(n109), .Z(n1140) );
  CENXL U1639 ( .A(n1735), .B(n109), .Z(n1143) );
  CND2IXL U1640 ( .B(n1736), .A(n109), .Z(n1144) );
  CENXL U1641 ( .A(n1680), .B(n109), .Z(n1142) );
  CENXL U1642 ( .A(n1681), .B(n109), .Z(n1141) );
  CENXL U1643 ( .A(a[28]), .B(n109), .Z(n1652) );
  CIVXL U1644 ( .A(n1698), .Z(n1473) );
  CND2IXL U1645 ( .B(n1736), .A(n1698), .Z(n1184) );
  CIVX3 U1646 ( .A(n48), .Z(n1731) );
  CENXL U1647 ( .A(n1716), .B(n152), .Z(n1341) );
  CIVXL U1648 ( .A(n339), .Z(n338) );
  CIVXL U1649 ( .A(n1696), .Z(n1475) );
  CND2IXL U1650 ( .B(n1736), .A(n1696), .Z(n1216) );
  CENXL U1651 ( .A(n1696), .B(n1692), .Z(n1202) );
  CENXL U1652 ( .A(n1696), .B(n1693), .Z(n1201) );
  CENXL U1653 ( .A(n1696), .B(n1690), .Z(n1204) );
  CENXL U1654 ( .A(n1696), .B(n1682), .Z(n1212) );
  CENXL U1655 ( .A(n1696), .B(n1683), .Z(n1211) );
  CENXL U1656 ( .A(n1696), .B(n1680), .Z(n1214) );
  CIVX1 U1657 ( .A(n912), .Z(n1620) );
  CIVX2 U1658 ( .A(n1620), .Z(n1621) );
  CIVX1 U1659 ( .A(n995), .Z(n1622) );
  CIVX2 U1660 ( .A(n1622), .Z(n1623) );
  CIVX1 U1661 ( .A(n996), .Z(n1624) );
  CIVX2 U1662 ( .A(n1624), .Z(n1625) );
  COND2XL U1663 ( .A(n91), .B(n1173), .C(n1172), .D(n89), .Z(n896) );
  COND2XL U1664 ( .A(n91), .B(n1176), .C(n1175), .D(n89), .Z(n899) );
  COND2XL U1665 ( .A(n91), .B(n1175), .C(n1174), .D(n89), .Z(n898) );
  COND2XL U1666 ( .A(n91), .B(n1174), .C(n1173), .D(n89), .Z(n897) );
  CFA1XL U1667 ( .A(n1047), .B(n1101), .CI(n1131), .CO(n840), .S(n841) );
  COND1X1 U1668 ( .A(n226), .B(n218), .C(n219), .Z(n217) );
  CIVX2 U1669 ( .A(n1565), .Z(n1626) );
  CIVX1 U1670 ( .A(n1565), .Z(n1627) );
  COND2XL U1671 ( .A(n102), .B(n1153), .C(n100), .D(n1152), .Z(n878) );
  COND2XL U1672 ( .A(n102), .B(n1154), .C(n100), .D(n1153), .Z(n879) );
  COND2XL U1673 ( .A(n102), .B(n1157), .C(n100), .D(n1156), .Z(n882) );
  COND2XL U1674 ( .A(n1159), .B(n102), .C(n100), .D(n1158), .Z(n884) );
  COND2XL U1675 ( .A(n85), .B(n1186), .C(n1185), .D(n1566), .Z(n908) );
  COND2XL U1676 ( .A(n85), .B(n1188), .C(n1187), .D(n1566), .Z(n910) );
  COND2XL U1677 ( .A(n85), .B(n1187), .C(n1186), .D(n1566), .Z(n909) );
  COND2XL U1678 ( .A(n85), .B(n1474), .C(n1627), .D(n1199), .Z(n856) );
  CND2X2 U1679 ( .A(n1449), .B(n1626), .Z(n85) );
  CIVX2 U1680 ( .A(a[0]), .Z(n1628) );
  CIVX1 U1681 ( .A(n1046), .Z(n1629) );
  CIVX2 U1682 ( .A(n1629), .Z(n1630) );
  CNIVX3 U1683 ( .A(n1702), .Z(n1632) );
  CFA1X1 U1684 ( .A(n1618), .B(n1054), .CI(n982), .CO(n578), .S(n579) );
  COND2X1 U1685 ( .A(n53), .B(n1264), .C(n1263), .D(n50), .Z(n982) );
  CIVX1 U1686 ( .A(a[14]), .Z(n1633) );
  CENXL U1687 ( .A(a[16]), .B(n1696), .Z(n1651) );
  CENXL U1688 ( .A(n1697), .B(n1680), .Z(n1197) );
  CANR1X1 U1689 ( .A(n1656), .B(n321), .C(n316), .Z(n314) );
  CIVXL U1690 ( .A(n1572), .Z(n278) );
  COND2XL U1691 ( .A(n44), .B(n1303), .C(n1302), .D(n42), .Z(n1020) );
  COND2XL U1692 ( .A(n44), .B(n1282), .C(n1281), .D(n42), .Z(n999) );
  CIVX4 U1693 ( .A(n1731), .Z(n1730) );
  COND2XL U1694 ( .A(n44), .B(n1283), .C(n1282), .D(n42), .Z(n1000) );
  CND2IXL U1695 ( .B(n1736), .A(n1714), .Z(n1360) );
  CNR2IXL U1696 ( .B(n1736), .A(n1649), .Z(n1075) );
  CND2X1 U1697 ( .A(n1637), .B(a[4]), .Z(n1639) );
  CIVXL U1698 ( .A(a[4]), .Z(n1638) );
  COND2XL U1699 ( .A(n27), .B(n1340), .C(n1649), .D(n1339), .Z(n1055) );
  COND2XL U1700 ( .A(n27), .B(n1342), .C(n1649), .D(n1341), .Z(n1057) );
  COND2XL U1701 ( .A(n27), .B(n1717), .C(n1360), .D(n1649), .Z(n863) );
  COND2XL U1702 ( .A(n27), .B(n1350), .C(n1649), .D(n1349), .Z(n1065) );
  COND2XL U1703 ( .A(n27), .B(n1341), .C(n1649), .D(n1340), .Z(n1056) );
  COND2XL U1704 ( .A(n27), .B(n1336), .C(n1649), .D(n1335), .Z(n1051) );
  COND2XL U1705 ( .A(n27), .B(n1335), .C(n1649), .D(n1334), .Z(n1050) );
  COND2XL U1706 ( .A(n27), .B(n1358), .C(n1649), .D(n1357), .Z(n1073) );
  COND2XL U1707 ( .A(n27), .B(n1333), .C(n1649), .D(n1332), .Z(n1048) );
  COND2XL U1708 ( .A(n27), .B(n1344), .C(n1649), .D(n1343), .Z(n1059) );
  COND2XL U1709 ( .A(n27), .B(n1351), .C(n1649), .D(n1350), .Z(n1066) );
  COND2XL U1710 ( .A(n27), .B(n1355), .C(n1649), .D(n1354), .Z(n1070) );
  COND2XL U1711 ( .A(n27), .B(n1353), .C(n1649), .D(n1352), .Z(n1068) );
  COND2XL U1712 ( .A(n27), .B(n1359), .C(n1649), .D(n1358), .Z(n1074) );
  COND2XL U1713 ( .A(n27), .B(n1354), .C(n1649), .D(n1353), .Z(n1069) );
  COND2XL U1714 ( .A(n27), .B(n1356), .C(n1649), .D(n1355), .Z(n1071) );
  COND2XL U1715 ( .A(n27), .B(n1334), .C(n1649), .D(n1333), .Z(n1049) );
  CND2XL U1716 ( .A(n1657), .B(n1659), .Z(n280) );
  CEOXL U1717 ( .A(n1080), .B(n1110), .Z(n1641) );
  CENX1 U1718 ( .A(n1730), .B(n1691), .Z(n1266) );
  CENX1 U1719 ( .A(n1730), .B(n1693), .Z(n1264) );
  CENX1 U1720 ( .A(n1730), .B(n1694), .Z(n1263) );
  CENX1 U1721 ( .A(n1730), .B(n150), .Z(n1262) );
  CEOX1 U1722 ( .A(n1641), .B(n980), .Z(n529) );
  CND2XL U1723 ( .A(n980), .B(n1110), .Z(n1642) );
  CND2XL U1724 ( .A(n980), .B(n1080), .Z(n1643) );
  CND2XL U1725 ( .A(n1110), .B(n1080), .Z(n1644) );
  CND3X1 U1726 ( .A(n1642), .B(n1643), .C(n1644), .Z(n528) );
  CNR2XL U1727 ( .A(n1261), .B(n50), .Z(n1646) );
  COR2X1 U1728 ( .A(n1645), .B(n1646), .Z(n980) );
  COND2XL U1729 ( .A(n9), .B(n1397), .C(n1564), .D(n1396), .Z(n1110) );
  CENX1 U1730 ( .A(n1730), .B(n151), .Z(n1261) );
  CIVX8 U1731 ( .A(n1731), .Z(n1729) );
  CNIVX1 U1732 ( .A(n144), .Z(n1692) );
  COND2XL U1733 ( .A(n18), .B(n1389), .C(n1670), .D(n1388), .Z(n1103) );
  CANR1X1 U1734 ( .A(n373), .B(n1664), .C(n370), .Z(n368) );
  CNR2IX1 U1735 ( .B(n1736), .A(n95), .Z(n895) );
  CANR1X1 U1736 ( .A(n331), .B(n339), .C(n332), .Z(n330) );
  CIVX2 U1737 ( .A(n3), .Z(n1704) );
  CND2XL U1738 ( .A(n1568), .B(n235), .Z(n171) );
  CND2X1 U1739 ( .A(n801), .B(n810), .Z(n337) );
  CND2XL U1740 ( .A(n412), .B(n375), .Z(n194) );
  COR2X1 U1741 ( .A(n1135), .B(n1105), .Z(n1665) );
  CEO3X1 U1742 ( .A(n434), .B(n416), .C(n432), .Z(n415) );
  CEO3X1 U1743 ( .A(n436), .B(n418), .C(n417), .Z(n416) );
  CEO3X1 U1744 ( .A(n422), .B(n421), .C(n440), .Z(n418) );
  CEO3X1 U1745 ( .A(n420), .B(n438), .C(n419), .Z(n417) );
  CEO3X1 U1746 ( .A(n452), .B(n450), .C(n448), .Z(n422) );
  COND2X1 U1747 ( .A(n69), .B(n1224), .C(n1223), .D(n66), .Z(n944) );
  CIVX1 U1748 ( .A(n1704), .Z(n1703) );
  COND2X1 U1749 ( .A(n91), .B(n1182), .C(n1181), .D(n89), .Z(n905) );
  CENX1 U1750 ( .A(n1721), .B(n151), .Z(n1313) );
  CNIVX3 U1751 ( .A(n134), .Z(n1687) );
  CEOXL U1752 ( .A(n236), .B(n171), .Z(product[26]) );
  CEOXL U1753 ( .A(n170), .B(n227), .Z(product[27]) );
  CND2XL U1754 ( .A(n388), .B(n226), .Z(n170) );
  CEOXL U1755 ( .A(n220), .B(n169), .Z(product[28]) );
  CAOR1X1 U1756 ( .A(n1654), .B(n213), .C(n210), .Z(n1647) );
  COND1X2 U1757 ( .A(n240), .B(n234), .C(n235), .Z(n229) );
  CND2XL U1758 ( .A(n390), .B(n240), .Z(n172) );
  CANR1X1 U1759 ( .A(n312), .B(n293), .C(n294), .Z(n292) );
  CNR2XL U1760 ( .A(n295), .B(n298), .Z(n293) );
  CND2XL U1761 ( .A(n1656), .B(n318), .Z(n182) );
  CANR1X1 U1762 ( .A(n308), .B(n1658), .C(n301), .Z(n299) );
  CIVX1 U1763 ( .A(n303), .Z(n301) );
  CEOXL U1764 ( .A(n177), .B(n286), .Z(product[20]) );
  CND2XL U1765 ( .A(n1657), .B(n285), .Z(n177) );
  CEOXL U1766 ( .A(n176), .B(n278), .Z(product[21]) );
  CEOXL U1767 ( .A(n181), .B(n1562), .Z(product[16]) );
  CND2XL U1768 ( .A(n399), .B(n306), .Z(n181) );
  CND2XL U1769 ( .A(n1659), .B(n290), .Z(n178) );
  CND2XL U1770 ( .A(n1658), .B(n303), .Z(n180) );
  CND2XL U1771 ( .A(n431), .B(n458), .Z(n207) );
  CND2XL U1772 ( .A(n1658), .B(n399), .Z(n298) );
  CNR2XL U1773 ( .A(n333), .B(n336), .Z(n331) );
  CNR2XL U1774 ( .A(n322), .B(n327), .Z(n320) );
  CND2XL U1775 ( .A(n1661), .B(n345), .Z(n187) );
  CND2XL U1776 ( .A(n1660), .B(n350), .Z(n188) );
  CND2XL U1777 ( .A(n402), .B(n328), .Z(n184) );
  CND2XL U1778 ( .A(n1662), .B(n356), .Z(n189) );
  CND2XL U1779 ( .A(n767), .B(n778), .Z(n323) );
  CND2XL U1780 ( .A(n430), .B(n415), .Z(n198) );
  CND2IXL U1781 ( .B(n358), .A(n359), .Z(n190) );
  CND2XL U1782 ( .A(n1666), .B(n364), .Z(n191) );
  CND2XL U1783 ( .A(n791), .B(n800), .Z(n334) );
  CND2IXL U1784 ( .B(n366), .A(n367), .Z(n192) );
  CND2XL U1785 ( .A(n1665), .B(n380), .Z(n195) );
  CEOXL U1786 ( .A(n376), .B(n194), .Z(product[3]) );
  CND2XL U1787 ( .A(n849), .B(n864), .Z(n375) );
  CAN2XL U1788 ( .A(n1569), .B(n383), .Z(product[1]) );
  CNR2IXL U1789 ( .B(n1736), .A(n114), .Z(n867) );
  CNR2IXL U1790 ( .B(n1736), .A(n89), .Z(n907) );
  CNR2IXL U1791 ( .B(n1736), .A(n100), .Z(n885) );
  COND2XL U1792 ( .A(n91), .B(n1180), .C(n1179), .D(n89), .Z(n903) );
  COND2XL U1793 ( .A(n97), .B(n1162), .C(n1161), .D(n95), .Z(n886) );
  COND2XL U1794 ( .A(n1138), .B(n115), .C(n114), .D(n1137), .Z(n866) );
  CNR2IXL U1795 ( .B(n1736), .A(n1564), .Z(product[0]) );
  COR2X2 U1796 ( .A(n1648), .B(n1669), .Z(n18) );
  CENX2 U1797 ( .A(n1697), .B(a[20]), .Z(n89) );
  CENXL U1798 ( .A(n1715), .B(a[6]), .Z(n33) );
  CENXL U1799 ( .A(n1631), .B(n156), .Z(n1401) );
  CNIVX2 U1800 ( .A(n104), .Z(n1701) );
  CND2IX1 U1801 ( .B(n1652), .A(n110), .Z(n112) );
  CND2XL U1802 ( .A(n1443), .B(n114), .Z(n115) );
  CNIVX4 U1803 ( .A(n140), .Z(n1690) );
  CIVX2 U1804 ( .A(n12), .Z(n1711) );
  CIVXL U1805 ( .A(n109), .Z(n1469) );
  CNR2X1 U1806 ( .A(n1571), .B(n239), .Z(n228) );
  COND1XL U1807 ( .A(n261), .B(n278), .C(n262), .Z(n260) );
  CND2XL U1808 ( .A(n391), .B(n250), .Z(n173) );
  COND1XL U1809 ( .A(n252), .B(n278), .C(n253), .Z(n251) );
  CENX1 U1810 ( .A(n241), .B(n172), .Z(product[25]) );
  COND1XL U1811 ( .A(n223), .B(n231), .C(n226), .Z(n222) );
  CANR1XL U1812 ( .A(n390), .B(n241), .C(n238), .Z(n236) );
  CANR1XL U1813 ( .A(n221), .B(n241), .C(n222), .Z(n220) );
  CNR2IXL U1814 ( .B(n228), .A(n223), .Z(n221) );
  CAN2X1 U1815 ( .A(n385), .B(n1654), .Z(n1653) );
  COND1XL U1816 ( .A(n295), .B(n299), .C(n296), .Z(n294) );
  CND2X1 U1817 ( .A(n320), .B(n1656), .Z(n313) );
  CNR2X1 U1818 ( .A(n563), .B(n586), .Z(n239) );
  CND2X1 U1819 ( .A(n397), .B(n296), .Z(n179) );
  CND2XL U1820 ( .A(n1567), .B(n270), .Z(n175) );
  COND1XL U1821 ( .A(n272), .B(n278), .C(n273), .Z(n271) );
  COND1XL U1822 ( .A(n305), .B(n1562), .C(n306), .Z(n304) );
  CENX1 U1823 ( .A(n291), .B(n178), .Z(product[19]) );
  CNR2X2 U1824 ( .A(n539), .B(n562), .Z(n234) );
  CANR1XL U1825 ( .A(n1659), .B(n291), .C(n288), .Z(n286) );
  CEOX1 U1826 ( .A(n183), .B(n324), .Z(product[14]) );
  CND2X1 U1827 ( .A(n401), .B(n323), .Z(n183) );
  CANR1XL U1828 ( .A(n402), .B(n329), .C(n326), .Z(n324) );
  CEOX1 U1829 ( .A(n182), .B(n319), .Z(product[15]) );
  CND2XL U1830 ( .A(n394), .B(n273), .Z(n176) );
  COR2X1 U1831 ( .A(n459), .B(n486), .Z(n1654) );
  CND2X1 U1832 ( .A(n513), .B(n538), .Z(n226) );
  CND2X1 U1833 ( .A(n609), .B(n630), .Z(n259) );
  COR2X1 U1834 ( .A(n609), .B(n630), .Z(n1655) );
  CND2X1 U1835 ( .A(n1661), .B(n1660), .Z(n340) );
  COND1XL U1836 ( .A(n337), .B(n333), .C(n334), .Z(n332) );
  CENX1 U1837 ( .A(n335), .B(n185), .Z(product[12]) );
  CND2X1 U1838 ( .A(n403), .B(n334), .Z(n185) );
  COND1XL U1839 ( .A(n336), .B(n338), .C(n337), .Z(n335) );
  CENX1 U1840 ( .A(n329), .B(n184), .Z(product[13]) );
  CNR2X1 U1841 ( .A(n767), .B(n778), .Z(n322) );
  CNR2X1 U1842 ( .A(n651), .B(n670), .Z(n272) );
  CNR2X1 U1843 ( .A(n739), .B(n752), .Z(n305) );
  COR2X1 U1844 ( .A(n753), .B(n766), .Z(n1656) );
  CEOX1 U1845 ( .A(n346), .B(n187), .Z(product[10]) );
  CANR1XL U1846 ( .A(n1660), .B(n351), .C(n348), .Z(n346) );
  CEOX1 U1847 ( .A(n186), .B(n338), .Z(product[11]) );
  CND2X1 U1848 ( .A(n404), .B(n337), .Z(n186) );
  COR2X1 U1849 ( .A(n671), .B(n688), .Z(n1657) );
  COR2X1 U1850 ( .A(n723), .B(n738), .Z(n1658) );
  COR2X1 U1851 ( .A(n689), .B(n706), .Z(n1659) );
  CND2X1 U1852 ( .A(n739), .B(n752), .Z(n306) );
  CND2X1 U1853 ( .A(n707), .B(n722), .Z(n296) );
  CND2X1 U1854 ( .A(n689), .B(n706), .Z(n290) );
  CND2X1 U1855 ( .A(n671), .B(n688), .Z(n285) );
  CND2X1 U1856 ( .A(n723), .B(n738), .Z(n303) );
  CND2X1 U1857 ( .A(n753), .B(n766), .Z(n318) );
  CENX1 U1858 ( .A(n189), .B(n357), .Z(product[8]) );
  COND1XL U1859 ( .A(n376), .B(n374), .C(n375), .Z(n373) );
  COND1XL U1860 ( .A(n368), .B(n366), .C(n367), .Z(n365) );
  CNR2X1 U1861 ( .A(n801), .B(n810), .Z(n336) );
  CNR2X1 U1862 ( .A(n791), .B(n800), .Z(n333) );
  CNR2X1 U1863 ( .A(n779), .B(n790), .Z(n327) );
  CND2X1 U1864 ( .A(n779), .B(n790), .Z(n328) );
  COR2X1 U1865 ( .A(n819), .B(n826), .Z(n1660) );
  COR2X1 U1866 ( .A(n811), .B(n818), .Z(n1661) );
  CND2X1 U1867 ( .A(n819), .B(n826), .Z(n350) );
  CND2X1 U1868 ( .A(n827), .B(n832), .Z(n356) );
  CND2X1 U1869 ( .A(n811), .B(n818), .Z(n345) );
  COR2X1 U1870 ( .A(n827), .B(n832), .Z(n1662) );
  COR2X1 U1871 ( .A(n430), .B(n415), .Z(n1663) );
  CENX1 U1872 ( .A(n193), .B(n373), .Z(product[4]) );
  CND2X1 U1873 ( .A(n1664), .B(n372), .Z(n193) );
  CENX1 U1874 ( .A(n195), .B(n381), .Z(product[2]) );
  CNR2X1 U1875 ( .A(n833), .B(n838), .Z(n358) );
  CNR2X1 U1876 ( .A(n849), .B(n864), .Z(n374) );
  CNR2X1 U1877 ( .A(n843), .B(n846), .Z(n366) );
  COR2X1 U1878 ( .A(n847), .B(n848), .Z(n1664) );
  CND2X1 U1879 ( .A(n833), .B(n838), .Z(n359) );
  CND2X1 U1880 ( .A(n1135), .B(n1105), .Z(n380) );
  CND2X1 U1881 ( .A(n847), .B(n848), .Z(n372) );
  CND2X1 U1882 ( .A(n839), .B(n842), .Z(n364) );
  CND2X1 U1883 ( .A(n843), .B(n846), .Z(n367) );
  COR2X1 U1884 ( .A(n839), .B(n842), .Z(n1666) );
  CENX1 U1885 ( .A(n1725), .B(n1690), .Z(n1292) );
  CENX1 U1886 ( .A(n1729), .B(n1692), .Z(n1265) );
  CENX1 U1887 ( .A(n1720), .B(n1689), .Z(n1320) );
  CENX1 U1888 ( .A(n1720), .B(n1688), .Z(n1321) );
  CENX1 U1889 ( .A(n1715), .B(n1687), .Z(n1351) );
  CENX1 U1890 ( .A(n1715), .B(n1688), .Z(n1350) );
  CENX1 U1891 ( .A(n1715), .B(n1689), .Z(n1349) );
  CENX1 U1892 ( .A(n1720), .B(n1690), .Z(n1319) );
  CENX1 U1893 ( .A(n1729), .B(n1685), .Z(n1272) );
  CENX1 U1894 ( .A(n1729), .B(n1687), .Z(n1270) );
  CENX1 U1895 ( .A(n1720), .B(n1691), .Z(n1318) );
  CENX1 U1896 ( .A(n1729), .B(n1684), .Z(n1273) );
  CENX1 U1897 ( .A(n1714), .B(n1692), .Z(n1346) );
  CENX1 U1898 ( .A(n1697), .B(n1692), .Z(n1185) );
  CENX1 U1899 ( .A(n1735), .B(n1631), .Z(n1423) );
  CENX1 U1900 ( .A(n1729), .B(n1686), .Z(n1271) );
  CENX1 U1901 ( .A(n1729), .B(n1680), .Z(n1277) );
  CENX1 U1902 ( .A(n1718), .B(n1681), .Z(n1328) );
  CENX1 U1903 ( .A(n1718), .B(n1682), .Z(n1327) );
  CENX1 U1904 ( .A(n1729), .B(n1683), .Z(n1274) );
  CENX1 U1905 ( .A(n1729), .B(n1681), .Z(n1276) );
  CENX1 U1906 ( .A(n1719), .B(n1686), .Z(n1323) );
  CENX1 U1907 ( .A(n1719), .B(n1685), .Z(n1324) );
  CENX1 U1908 ( .A(n1718), .B(n1683), .Z(n1326) );
  CENX1 U1909 ( .A(n1729), .B(n1682), .Z(n1275) );
  CENX1 U1910 ( .A(n1707), .B(n1682), .Z(n1387) );
  CENX1 U1911 ( .A(n1707), .B(n1683), .Z(n1386) );
  CENX1 U1912 ( .A(n1708), .B(n1687), .Z(n1382) );
  CENX1 U1913 ( .A(n1709), .B(n1694), .Z(n1375) );
  CENX1 U1914 ( .A(n1706), .B(n1685), .Z(n1384) );
  CENX1 U1915 ( .A(n1707), .B(n1684), .Z(n1385) );
  CENX1 U1916 ( .A(n1706), .B(n1686), .Z(n1383) );
  CNR2IXL U1917 ( .B(n1736), .A(n1670), .Z(n1105) );
  CENX1 U1918 ( .A(n1697), .B(n1685), .Z(n1192) );
  CENX1 U1919 ( .A(n1697), .B(n1686), .Z(n1191) );
  CENX1 U1920 ( .A(n1697), .B(n1684), .Z(n1193) );
  CENX1 U1921 ( .A(n1730), .B(n1690), .Z(n1267) );
  CENX1 U1922 ( .A(n1697), .B(n1682), .Z(n1195) );
  CENX1 U1923 ( .A(n1726), .B(n1694), .Z(n1288) );
  CENX1 U1924 ( .A(n1725), .B(n1689), .Z(n1293) );
  CENX1 U1925 ( .A(n1724), .B(n1688), .Z(n1294) );
  CENX1 U1926 ( .A(n1724), .B(n1687), .Z(n1295) );
  CENX1 U1927 ( .A(n1725), .B(n1692), .Z(n1290) );
  CENX1 U1928 ( .A(n1726), .B(n1693), .Z(n1289) );
  CENX1 U1929 ( .A(n1724), .B(n1685), .Z(n1297) );
  CENX1 U1930 ( .A(n1724), .B(n1684), .Z(n1298) );
  CENX1 U1931 ( .A(n1724), .B(n1683), .Z(n1299) );
  CENX1 U1932 ( .A(n1724), .B(n1681), .Z(n1301) );
  CENX1 U1933 ( .A(n1724), .B(n1680), .Z(n1302) );
  CENX1 U1934 ( .A(n1697), .B(n1691), .Z(n1186) );
  CENX1 U1935 ( .A(n1697), .B(n1690), .Z(n1187) );
  CENX1 U1936 ( .A(n1697), .B(n1687), .Z(n1190) );
  CENX1 U1937 ( .A(n1697), .B(n1688), .Z(n1189) );
  CENX1 U1938 ( .A(n1714), .B(n1681), .Z(n1357) );
  CENX1 U1939 ( .A(n1714), .B(n1680), .Z(n1358) );
  CENX1 U1940 ( .A(n1631), .B(n1694), .Z(n1408) );
  CENX1 U1941 ( .A(n1632), .B(n1693), .Z(n1409) );
  CENX1 U1942 ( .A(n1631), .B(n1680), .Z(n1422) );
  CENX1 U1943 ( .A(n1631), .B(n1681), .Z(n1421) );
  CENX1 U1944 ( .A(n1631), .B(n1683), .Z(n1419) );
  CENX1 U1945 ( .A(n1632), .B(n1684), .Z(n1418) );
  CENX1 U1946 ( .A(n1632), .B(n1687), .Z(n1415) );
  CENX1 U1947 ( .A(n1713), .B(n1683), .Z(n1355) );
  CENX1 U1948 ( .A(n1631), .B(n1685), .Z(n1417) );
  CENX1 U1949 ( .A(n1632), .B(n1686), .Z(n1416) );
  CENX1 U1950 ( .A(n1632), .B(n1690), .Z(n1412) );
  CENX1 U1951 ( .A(n1713), .B(n1686), .Z(n1352) );
  CENX1 U1952 ( .A(n1631), .B(n1692), .Z(n1410) );
  CENX1 U1953 ( .A(n1632), .B(n1691), .Z(n1411) );
  CENX1 U1954 ( .A(n1713), .B(n1685), .Z(n1353) );
  CENX1 U1955 ( .A(n1713), .B(n1684), .Z(n1354) );
  CENX1 U1956 ( .A(n1632), .B(n1689), .Z(n1413) );
  CENX1 U1957 ( .A(n1632), .B(n1688), .Z(n1414) );
  CENX1 U1958 ( .A(n1730), .B(n1688), .Z(n1269) );
  CENX1 U1959 ( .A(n1733), .B(n1692), .Z(n1242) );
  CENX1 U1960 ( .A(n1732), .B(n1686), .Z(n1248) );
  CENX1 U1961 ( .A(n1730), .B(n1689), .Z(n1268) );
  CENX1 U1962 ( .A(n1718), .B(n1687), .Z(n1322) );
  CENX1 U1963 ( .A(n1735), .B(n1697), .Z(n1198) );
  CENX1 U1964 ( .A(n1732), .B(n1687), .Z(n1247) );
  CENX1 U1965 ( .A(n1732), .B(n1683), .Z(n1251) );
  CENX1 U1966 ( .A(n1733), .B(n1693), .Z(n1241) );
  CENX1 U1967 ( .A(n1733), .B(n1694), .Z(n1240) );
  CENX1 U1968 ( .A(n1718), .B(n1680), .Z(n1329) );
  CENX1 U1969 ( .A(n1637), .B(n1680), .Z(n1389) );
  CENX1 U1970 ( .A(n1637), .B(n1690), .Z(n1379) );
  CENX1 U1971 ( .A(n1735), .B(n1710), .Z(n1390) );
  CENX1 U1972 ( .A(n1735), .B(n1721), .Z(n1330) );
  CENX1 U1973 ( .A(n1735), .B(n1730), .Z(n1278) );
  CENX1 U1974 ( .A(n1736), .B(n1733), .Z(n1255) );
  CNR2IX1 U1975 ( .B(n1736), .A(n42), .Z(n1021) );
  CEOX1 U1976 ( .A(n872), .B(n886), .Z(n429) );
  CENX1 U1977 ( .A(n1718), .B(b[25]), .Z(n1305) );
  CENX1 U1978 ( .A(n1729), .B(n155), .Z(n1257) );
  CENX1 U1979 ( .A(n1637), .B(b[29]), .Z(n1361) );
  CENX1 U1980 ( .A(n1733), .B(n153), .Z(n1236) );
  CENX1 U1981 ( .A(n1719), .B(n154), .Z(n1310) );
  CENX1 U1982 ( .A(n1723), .B(n155), .Z(n1282) );
  CENX1 U1983 ( .A(n1710), .B(n151), .Z(n1373) );
  CENX1 U1984 ( .A(n1712), .B(n157), .Z(n1336) );
  CENX1 U1985 ( .A(n1716), .B(n151), .Z(n1342) );
  CENX1 U1986 ( .A(n1719), .B(n155), .Z(n1309) );
  CENX1 U1987 ( .A(n1718), .B(n150), .Z(n1314) );
  CENX1 U1988 ( .A(n1710), .B(n150), .Z(n1374) );
  CENX1 U1989 ( .A(n109), .B(a[30]), .Z(n114) );
  CENX1 U1990 ( .A(n1705), .B(b[24]), .Z(n1366) );
  CENX1 U1991 ( .A(n1631), .B(b[31]), .Z(n1392) );
  CENX1 U1992 ( .A(n1714), .B(b[27]), .Z(n1332) );
  CENX1 U1993 ( .A(n1729), .B(n153), .Z(n1259) );
  CENX1 U1994 ( .A(n1705), .B(b[25]), .Z(n1365) );
  CENX1 U1995 ( .A(n1723), .B(n154), .Z(n1283) );
  CENX1 U1996 ( .A(n1723), .B(n153), .Z(n1284) );
  CENX1 U1997 ( .A(n1723), .B(n156), .Z(n1281) );
  CENXL U1998 ( .A(n1631), .B(n157), .Z(n1400) );
  CENX1 U1999 ( .A(n1632), .B(n151), .Z(n1406) );
  CENX1 U2000 ( .A(n1714), .B(n153), .Z(n1340) );
  CENX1 U2001 ( .A(n1631), .B(b[24]), .Z(n1399) );
  CENX1 U2002 ( .A(n1632), .B(n154), .Z(n1403) );
  CENX1 U2003 ( .A(n1631), .B(n150), .Z(n1407) );
  CENX1 U2004 ( .A(n1632), .B(b[26]), .Z(n1397) );
  CENX1 U2005 ( .A(n1631), .B(b[27]), .Z(n1396) );
  CENX1 U2006 ( .A(n1632), .B(b[25]), .Z(n1398) );
  CENX1 U2007 ( .A(n1716), .B(b[24]), .Z(n1335) );
  CENX1 U2008 ( .A(n1632), .B(b[28]), .Z(n1395) );
  CENX1 U2009 ( .A(n1712), .B(b[25]), .Z(n1334) );
  CENX1 U2010 ( .A(n1632), .B(b[30]), .Z(n1393) );
  CENX1 U2011 ( .A(n1715), .B(b[26]), .Z(n1333) );
  CENX1 U2012 ( .A(n1631), .B(b[29]), .Z(n1394) );
  CND2X2 U2013 ( .A(n1455), .B(n1673), .Z(n36) );
  CENX1 U2014 ( .A(n1680), .B(n113), .Z(n1137) );
  CENX1 U2015 ( .A(n1735), .B(n113), .Z(n1138) );
  CENX1 U2016 ( .A(n1718), .B(n156), .Z(n1308) );
  CENX1 U2017 ( .A(n1733), .B(n150), .Z(n1239) );
  CENX1 U2018 ( .A(n1718), .B(b[24]), .Z(n1306) );
  CENX1 U2019 ( .A(n1733), .B(n151), .Z(n1238) );
  CENX1 U2020 ( .A(n1718), .B(n157), .Z(n1307) );
  CENX1 U2021 ( .A(n1637), .B(b[26]), .Z(n1364) );
  CENX1 U2022 ( .A(n1708), .B(b[27]), .Z(n1363) );
  CENX1 U2023 ( .A(n1707), .B(b[28]), .Z(n1362) );
  CEOX1 U2024 ( .A(a[18]), .B(n1697), .Z(n1449) );
  CEOX2 U2025 ( .A(a[12]), .B(n1733), .Z(n1452) );
  CEOX2 U2026 ( .A(n1721), .B(a[8]), .Z(n1668) );
  CEOX1 U2027 ( .A(a[30]), .B(n113), .Z(n1443) );
  COND2XL U2028 ( .A(n69), .B(n1218), .C(n1217), .D(n66), .Z(n938) );
  COND2XL U2029 ( .A(n69), .B(n1219), .C(n1218), .D(n66), .Z(n939) );
  COND2XL U2030 ( .A(n69), .B(n1220), .C(n1219), .D(n66), .Z(n940) );
  COND2XL U2031 ( .A(n69), .B(n1221), .C(n1220), .D(n66), .Z(n941) );
  CNR2IXL U2032 ( .B(n1736), .A(n66), .Z(n955) );
  COND2XL U2033 ( .A(n69), .B(n1586), .C(n66), .D(n1235), .Z(n858) );
  COND2XL U2034 ( .A(n69), .B(n1230), .C(n1229), .D(n66), .Z(n950) );
  CIVX1 U2035 ( .A(n1671), .Z(n1672) );
  CND2X1 U2036 ( .A(n1136), .B(n865), .Z(n383) );
  COND2X1 U2037 ( .A(n61), .B(n1253), .C(n1252), .D(n58), .Z(n972) );
  CENX1 U2038 ( .A(n1715), .B(a[6]), .Z(n1673) );
  CIVX1 U2039 ( .A(n1717), .Z(n1715) );
  COND2X1 U2040 ( .A(n77), .B(n1214), .C(n1213), .D(n74), .Z(n935) );
  CIVX2 U2041 ( .A(n39), .Z(n1728) );
  CNR2X1 U2042 ( .A(n245), .B(n261), .Z(n243) );
  COND2XL U2043 ( .A(n77), .B(n1201), .C(n1200), .D(n74), .Z(n922) );
  COND2XL U2044 ( .A(n77), .B(n1203), .C(n1202), .D(n74), .Z(n924) );
  COND2XL U2045 ( .A(n77), .B(n1204), .C(n1203), .D(n74), .Z(n925) );
  COND2XL U2046 ( .A(n77), .B(n1202), .C(n1201), .D(n74), .Z(n923) );
  COND2XL U2047 ( .A(n1215), .B(n77), .C(n1214), .D(n74), .Z(n936) );
  CND2IXL U2048 ( .B(n1736), .A(n1695), .Z(n1235) );
  CEOXL U2049 ( .A(n368), .B(n192), .Z(product[5]) );
  CND2X1 U2050 ( .A(n487), .B(n512), .Z(n219) );
  CND2XL U2051 ( .A(n387), .B(n219), .Z(n169) );
  CND2X1 U2052 ( .A(n459), .B(n486), .Z(n212) );
  CND2XL U2053 ( .A(n1654), .B(n212), .Z(n168) );
  CIVXL U2054 ( .A(n1679), .Z(n1674) );
  CIVX1 U2055 ( .A(n1674), .Z(n1675) );
  CFA1XL U2056 ( .A(n955), .B(n993), .CI(n973), .CO(n776), .S(n777) );
  CFA1XL U2057 ( .A(n997), .B(n1043), .CI(n1019), .CO(n816), .S(n817) );
  COND2X1 U2058 ( .A(n36), .B(n1310), .C(n1309), .D(n1679), .Z(n1026) );
  COND2X1 U2059 ( .A(n61), .B(n1250), .C(n1249), .D(n58), .Z(n969) );
  CENX1 U2060 ( .A(n1714), .B(n1693), .Z(n1345) );
  CENX1 U2061 ( .A(n1714), .B(n1690), .Z(n1348) );
  CENX1 U2062 ( .A(n1714), .B(n1691), .Z(n1347) );
  COND1XL U2063 ( .A(n212), .B(n206), .C(n207), .Z(n1676) );
  COND2X1 U2064 ( .A(n36), .B(n1311), .C(n1310), .D(n1679), .Z(n1027) );
  CFA1X1 U2065 ( .A(n1030), .B(n629), .CI(n1114), .CO(n620), .S(n621) );
  COND2XL U2066 ( .A(n53), .B(n1258), .C(n1257), .D(n50), .Z(n976) );
  COND2XL U2067 ( .A(n53), .B(n1274), .C(n1273), .D(n50), .Z(n992) );
  CNR2IXL U2068 ( .B(n1736), .A(n50), .Z(n997) );
  COND2XL U2069 ( .A(n53), .B(n1260), .C(n1259), .D(n50), .Z(n978) );
  COND2XL U2070 ( .A(n53), .B(n1261), .C(n1260), .D(n50), .Z(n979) );
  COND2XL U2071 ( .A(n53), .B(n1278), .C(n1277), .D(n50), .Z(n996) );
  COND2XL U2072 ( .A(n53), .B(n1269), .C(n1268), .D(n50), .Z(n987) );
  COND2XL U2073 ( .A(n53), .B(n1271), .C(n1270), .D(n50), .Z(n989) );
  COND2XL U2074 ( .A(n53), .B(n1277), .C(n1276), .D(n50), .Z(n995) );
  COND2XL U2075 ( .A(n53), .B(n1276), .C(n1275), .D(n50), .Z(n994) );
  CENX1 U2076 ( .A(n188), .B(n351), .Z(product[9]) );
  COND2XL U2077 ( .A(n36), .B(n1306), .C(n1305), .D(n1675), .Z(n1022) );
  COND2XL U2078 ( .A(n36), .B(n1328), .C(n1327), .D(n1675), .Z(n1044) );
  COND2XL U2079 ( .A(n36), .B(n1307), .C(n1306), .D(n1675), .Z(n1023) );
  COND2XL U2080 ( .A(n36), .B(n1308), .C(n1307), .D(n1675), .Z(n1024) );
  COND2XL U2081 ( .A(n36), .B(n1326), .C(n1325), .D(n1675), .Z(n1042) );
  COND2XL U2082 ( .A(n36), .B(n1330), .C(n1329), .D(n1675), .Z(n1046) );
  COND2XL U2083 ( .A(n36), .B(n1722), .C(n1331), .D(n1675), .Z(n862) );
  COND2XL U2084 ( .A(n36), .B(n1323), .C(n1322), .D(n1679), .Z(n1039) );
  CNR2IXL U2085 ( .B(n1736), .A(n1679), .Z(n1047) );
  COND2XL U2086 ( .A(n36), .B(n1329), .C(n1328), .D(n1679), .Z(n1045) );
  COND2XL U2087 ( .A(n36), .B(n1309), .C(n1308), .D(n1679), .Z(n1025) );
  COND2XL U2088 ( .A(n36), .B(n1317), .C(n1316), .D(n1679), .Z(n1033) );
  COND2XL U2089 ( .A(n36), .B(n1324), .C(n1323), .D(n1679), .Z(n1040) );
  COND2XL U2090 ( .A(n36), .B(n1325), .C(n1324), .D(n1679), .Z(n1041) );
  COND2XL U2091 ( .A(n36), .B(n1319), .C(n1318), .D(n1679), .Z(n1035) );
  COND2XL U2092 ( .A(n36), .B(n1327), .C(n1326), .D(n1679), .Z(n1043) );
  CENX1 U2093 ( .A(n1631), .B(n155), .Z(n1402) );
  CIVX1 U2094 ( .A(n1717), .Z(n1713) );
  CIVX1 U2095 ( .A(n1582), .Z(n1727) );
  CENX1 U2096 ( .A(n1705), .B(n156), .Z(n1368) );
  COND2X1 U2097 ( .A(n18), .B(n1367), .C(n1670), .D(n1366), .Z(n1081) );
  COND2XL U2098 ( .A(n18), .B(n1362), .C(n1670), .D(n1361), .Z(n1076) );
  COND2XL U2099 ( .A(n18), .B(n1363), .C(n1670), .D(n1362), .Z(n1077) );
  COND2XL U2100 ( .A(n18), .B(n1711), .C(n1391), .D(n1670), .Z(n864) );
  COND2XL U2101 ( .A(n18), .B(n1388), .C(n1670), .D(n1387), .Z(n1102) );
  COND2XL U2102 ( .A(n18), .B(n1385), .C(n1670), .D(n1384), .Z(n1099) );
  COND2XL U2103 ( .A(n18), .B(n1383), .C(n1670), .D(n1382), .Z(n1097) );
  COND2XL U2104 ( .A(n18), .B(n1386), .C(n1670), .D(n1385), .Z(n1100) );
  COND2XL U2105 ( .A(n18), .B(n1384), .C(n1670), .D(n1383), .Z(n1098) );
  COND2XL U2106 ( .A(n18), .B(n1390), .C(n1670), .D(n1389), .Z(n1104) );
  COND2XL U2107 ( .A(n18), .B(n1365), .C(n1670), .D(n1364), .Z(n1079) );
  COND2XL U2108 ( .A(n18), .B(n1364), .C(n1670), .D(n1363), .Z(n1078) );
  COND2XL U2109 ( .A(n18), .B(n1370), .C(n1670), .D(n1369), .Z(n1084) );
  COND2XL U2110 ( .A(n18), .B(n1387), .C(n1670), .D(n1386), .Z(n1101) );
  COND2XL U2111 ( .A(n18), .B(n1379), .C(n1670), .D(n1378), .Z(n1093) );
  COND2XL U2112 ( .A(n18), .B(n1380), .C(n1670), .D(n1379), .Z(n1094) );
  COND2XL U2113 ( .A(n18), .B(n1382), .C(n1670), .D(n1381), .Z(n1096) );
  COND2XL U2114 ( .A(n18), .B(n1376), .C(n1670), .D(n1375), .Z(n1090) );
  COND2XL U2115 ( .A(n9), .B(n1704), .C(n1564), .D(n1424), .Z(n865) );
  COND2XL U2116 ( .A(n18), .B(n1366), .C(n1670), .D(n1365), .Z(n1080) );
  CENX1 U2117 ( .A(n1709), .B(n1693), .Z(n1376) );
  CENX1 U2118 ( .A(n1709), .B(n1691), .Z(n1378) );
  CENX1 U2119 ( .A(n1709), .B(n1692), .Z(n1377) );
  CANR1XL U2120 ( .A(n320), .B(n329), .C(n321), .Z(n319) );
  CENX1 U2121 ( .A(n1718), .B(n1684), .Z(n1325) );
  CENX1 U2122 ( .A(n1708), .B(n1688), .Z(n1381) );
  CENX1 U2123 ( .A(n1708), .B(n1689), .Z(n1380) );
  CND2XL U2124 ( .A(n1655), .B(n259), .Z(n174) );
  CND2XL U2125 ( .A(n263), .B(n1655), .Z(n252) );
  CANR1XL U2126 ( .A(n1655), .B(n264), .C(n257), .Z(n253) );
  CIVXL U2127 ( .A(n218), .Z(n387) );
  CNR2X2 U2128 ( .A(n487), .B(n512), .Z(n218) );
  CND2X1 U2129 ( .A(n216), .B(n228), .Z(n214) );
  CEOXL U2130 ( .A(n360), .B(n190), .Z(product[7]) );
  CENX1 U2131 ( .A(n1707), .B(n1681), .Z(n1388) );
  CENX1 U2132 ( .A(n1716), .B(n150), .Z(n1343) );
  COND2X1 U2133 ( .A(n18), .B(n1369), .C(n1670), .D(n1368), .Z(n1083) );
  CENX1 U2134 ( .A(n1724), .B(n1686), .Z(n1296) );
  CANR1X2 U2135 ( .A(n275), .B(n1567), .C(n268), .Z(n262) );
  COND2X1 U2136 ( .A(n61), .B(n1249), .C(n1248), .D(n58), .Z(n968) );
  COND2X1 U2137 ( .A(n36), .B(n1315), .C(n1314), .D(n1679), .Z(n1031) );
  CIVX1 U2138 ( .A(n965), .Z(n1677) );
  CIVX2 U2139 ( .A(n1677), .Z(n1678) );
  COND2XL U2140 ( .A(n61), .B(n1237), .C(n1236), .D(n58), .Z(n956) );
  COND2XL U2141 ( .A(n61), .B(n1238), .C(n1237), .D(n58), .Z(n957) );
  COND2XL U2142 ( .A(n61), .B(n1240), .C(n1239), .D(n58), .Z(n959) );
  COND2XL U2143 ( .A(n61), .B(n1251), .C(n1250), .D(n58), .Z(n970) );
  COND2XL U2144 ( .A(n53), .B(n1731), .C(n1279), .D(n50), .Z(n860) );
  COND2XL U2145 ( .A(n61), .B(n1239), .C(n1238), .D(n58), .Z(n958) );
  CNR2IXL U2146 ( .B(n1736), .A(n58), .Z(n975) );
  COND2XL U2147 ( .A(n61), .B(n1734), .C(n1256), .D(n58), .Z(n859) );
  COND2XL U2148 ( .A(n61), .B(n1245), .C(n1244), .D(n58), .Z(n964) );
  COND2XL U2149 ( .A(n61), .B(n1242), .C(n1241), .D(n58), .Z(n961) );
  COND2XL U2150 ( .A(n61), .B(n1255), .C(n1254), .D(n58), .Z(n974) );
  COND2XL U2151 ( .A(n61), .B(n1252), .C(n1251), .D(n58), .Z(n971) );
  COND2XL U2152 ( .A(n61), .B(n1241), .C(n1240), .D(n58), .Z(n960) );
  COND2XL U2153 ( .A(n61), .B(n1248), .C(n1247), .D(n58), .Z(n967) );
  COND2XL U2154 ( .A(n61), .B(n1246), .C(n1245), .D(n58), .Z(n965) );
  COND1XL U2155 ( .A(n298), .B(n1562), .C(n299), .Z(n297) );
  CENX1 U2156 ( .A(n1707), .B(n153), .Z(n1371) );
  COND2XL U2157 ( .A(n36), .B(n1314), .C(n1313), .D(n1679), .Z(n1030) );
  CENX1 U2158 ( .A(n1718), .B(n1693), .Z(n1316) );
  CENX1 U2159 ( .A(n1718), .B(n1694), .Z(n1315) );
  CENX1 U2160 ( .A(n1706), .B(n154), .Z(n1370) );
  CENX1 U2161 ( .A(n1724), .B(n1691), .Z(n1291) );
  CIVX1 U2162 ( .A(n1728), .Z(n1724) );
  CIVX1 U2163 ( .A(n1582), .Z(n1726) );
  CIVX2 U2164 ( .A(n1582), .Z(n1725) );
  CENX1 U2165 ( .A(n1726), .B(n151), .Z(n1286) );
  CENX1 U2166 ( .A(n1726), .B(n150), .Z(n1287) );
  CIVXL U2167 ( .A(n262), .Z(n264) );
  COND2X1 U2168 ( .A(n18), .B(n1368), .C(n1670), .D(n1367), .Z(n1082) );
  CENX1 U2169 ( .A(n1718), .B(n153), .Z(n1311) );
  CIVX2 U2170 ( .A(n1722), .Z(n1718) );
  CIVX2 U2171 ( .A(n30), .Z(n1722) );
  CIVX1 U2172 ( .A(n1711), .Z(n1710) );
  CNR2X1 U2173 ( .A(n218), .B(n223), .Z(n216) );
  CND2X4 U2174 ( .A(n1458), .B(n1564), .Z(n9) );
  CENX4 U2175 ( .A(n1729), .B(a[12]), .Z(n58) );
  CND2X4 U2176 ( .A(n1452), .B(n58), .Z(n61) );
  CENX4 U2177 ( .A(n1732), .B(n1634), .Z(n66) );
  CIVXL U2178 ( .A(n1711), .Z(n1705) );
  CIVXL U2179 ( .A(n1711), .Z(n1706) );
  CIVXL U2180 ( .A(n1711), .Z(n1708) );
  CIVXL U2181 ( .A(n1711), .Z(n1709) );
  CIVXL U2182 ( .A(n1717), .Z(n1712) );
  CIVXL U2183 ( .A(n1717), .Z(n1716) );
  CIVX2 U2184 ( .A(n21), .Z(n1717) );
  CIVXL U2185 ( .A(n1722), .Z(n1719) );
  CIVXL U2186 ( .A(n1722), .Z(n1720) );
  CIVXL U2187 ( .A(n1728), .Z(n1723) );
  CIVX2 U2188 ( .A(n374), .Z(n412) );
  CIVX2 U2189 ( .A(n336), .Z(n404) );
  CIVX2 U2190 ( .A(n333), .Z(n403) );
  CIVX2 U2191 ( .A(n295), .Z(n397) );
  CIVX2 U2192 ( .A(n223), .Z(n388) );
  CIVX2 U2193 ( .A(n383), .Z(n381) );
  CIVX2 U2194 ( .A(n380), .Z(n378) );
  CIVX2 U2195 ( .A(n372), .Z(n370) );
  CIVX2 U2196 ( .A(n364), .Z(n362) );
  CIVX2 U2197 ( .A(n356), .Z(n354) );
  CIVX2 U2198 ( .A(n350), .Z(n348) );
  CIVX2 U2199 ( .A(n345), .Z(n343) );
  CIVX2 U2200 ( .A(n328), .Z(n326) );
  CIVX2 U2201 ( .A(n327), .Z(n402) );
  CIVX2 U2202 ( .A(n318), .Z(n316) );
  CIVX2 U2203 ( .A(n306), .Z(n308) );
  CIVX2 U2204 ( .A(n305), .Z(n399) );
  CIVX2 U2205 ( .A(n290), .Z(n288) );
  CIVX2 U2206 ( .A(n285), .Z(n283) );
  CIVX2 U2207 ( .A(n273), .Z(n275) );
  CIVX2 U2208 ( .A(n270), .Z(n268) );
  CIVX2 U2209 ( .A(n249), .Z(n391) );
  CIVX2 U2210 ( .A(n240), .Z(n238) );
  CIVX2 U2211 ( .A(n212), .Z(n210) );
  CIVX2 U2212 ( .A(n1697), .Z(n1474) );
  CIVX2 U2213 ( .A(n1701), .Z(n1470) );
  CIVX2 U2214 ( .A(n113), .Z(n1468) );
endmodule


module calc_DW_mult_uns_18 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n3, n6, n9, n12, n15, n18, n21, n27, n30, n36, n39, n44, n48, n50,
         n53, n55, n58, n61, n63, n66, n69, n71, n74, n77, n79, n82, n85, n87,
         n89, n91, n93, n95, n97, n99, n100, n102, n104, n105, n107, n109,
         n110, n112, n113, n114, n115, n116, n120, n122, n124, n126, n128,
         n130, n132, n134, n136, n138, n140, n142, n144, n146, n148, n150,
         n151, n152, n153, n154, n155, n156, n157, n168, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n198, n199, n205, n207, n208, n210, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n226, n227, n228, n229,
         n234, n235, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n248, n250, n251, n252, n253, n257, n259, n260, n261, n262, n263,
         n264, n268, n270, n271, n272, n273, n275, n278, n279, n280, n281,
         n283, n285, n286, n288, n290, n292, n293, n294, n295, n296, n297,
         n298, n299, n301, n303, n304, n305, n306, n308, n311, n312, n313,
         n314, n316, n318, n319, n320, n321, n322, n323, n324, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n343, n345, n346, n348, n350, n351, n352, n354,
         n356, n357, n358, n359, n360, n362, n364, n365, n366, n367, n368,
         n370, n372, n373, n374, n375, n376, n378, n380, n381, n383, n387,
         n388, n389, n390, n394, n397, n399, n401, n402, n403, n404, n412,
         n415, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1443, n1445, n1447, n1448,
         n1449, n1450, n1451, n1452, n1455, n1457, n1458, n1468, n1469, n1470,
         n1472, n1473, n1474, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746;
  assign n3 = a[1];
  assign n12 = a[3];
  assign n21 = a[5];
  assign n30 = a[7];
  assign n39 = a[9];
  assign n48 = a[11];
  assign n55 = a[13];
  assign n63 = a[15];
  assign n71 = a[17];
  assign n79 = a[19];
  assign n87 = a[21];
  assign n93 = a[23];
  assign n99 = a[25];
  assign n104 = a[27];
  assign n109 = a[29];
  assign n113 = a[31];
  assign n116 = b[0];
  assign n120 = b[1];
  assign n122 = b[2];
  assign n124 = b[3];
  assign n126 = b[4];
  assign n128 = b[5];
  assign n130 = b[6];
  assign n132 = b[7];
  assign n134 = b[8];
  assign n136 = b[9];
  assign n138 = b[10];
  assign n140 = b[11];
  assign n142 = b[12];
  assign n144 = b[13];
  assign n146 = b[14];
  assign n148 = b[15];
  assign n150 = b[16];
  assign n151 = b[17];
  assign n152 = b[18];
  assign n153 = b[19];
  assign n154 = b[20];
  assign n155 = b[21];
  assign n156 = b[22];
  assign n157 = b[23];

  CEO3X2 U410 ( .A(n420), .B(n438), .C(n419), .Z(n417) );
  CEO3X2 U411 ( .A(n422), .B(n421), .C(n440), .Z(n418) );
  CEO3X2 U412 ( .A(n444), .B(n423), .C(n442), .Z(n419) );
  CEO3X2 U413 ( .A(n425), .B(n424), .C(n446), .Z(n420) );
  CEO3X2 U414 ( .A(n428), .B(n427), .C(n426), .Z(n421) );
  CEO3X2 U416 ( .A(n456), .B(n429), .C(n454), .Z(n423) );
  CEO3X2 U417 ( .A(n956), .B(n1022), .C(n1106), .Z(n424) );
  CEO3X2 U418 ( .A(n938), .B(n998), .C(n1076), .Z(n425) );
  CEO3X2 U419 ( .A(n866), .B(n976), .C(n1048), .Z(n426) );
  CEO3X2 U420 ( .A(n868), .B(n896), .C(n922), .Z(n427) );
  CEO3X2 U421 ( .A(n878), .B(n850), .C(n908), .Z(n428) );
  CFA1X1 U423 ( .A(n435), .B(n433), .CI(n460), .CO(n430), .S(n431) );
  CFA1X1 U424 ( .A(n439), .B(n462), .CI(n437), .CO(n432), .S(n433) );
  CFA1X1 U425 ( .A(n441), .B(n464), .CI(n466), .CO(n434), .S(n435) );
  CFA1X1 U426 ( .A(n445), .B(n443), .CI(n468), .CO(n436), .S(n437) );
  CFA1X1 U427 ( .A(n472), .B(n447), .CI(n470), .CO(n438), .S(n439) );
  CFA1X1 U428 ( .A(n474), .B(n449), .CI(n451), .CO(n440), .S(n441) );
  CFA1X1 U429 ( .A(n457), .B(n453), .CI(n455), .CO(n442), .S(n443) );
  CFA1X1 U430 ( .A(n480), .B(n476), .CI(n478), .CO(n444), .S(n445) );
  CFA1X1 U431 ( .A(n1023), .B(n482), .CI(n484), .CO(n446), .S(n447) );
  CFA1X1 U432 ( .A(n957), .B(n1077), .CI(n1107), .CO(n448), .S(n449) );
  CFA1X1 U433 ( .A(n939), .B(n1049), .CI(n999), .CO(n450), .S(n451) );
  CFA1X1 U435 ( .A(n869), .B(n1564), .CI(n887), .CO(n454), .S(n455) );
  CFA1X1 U436 ( .A(n867), .B(n873), .CI(n879), .CO(n456), .S(n457) );
  CFA1X1 U437 ( .A(n463), .B(n461), .CI(n488), .CO(n458), .S(n459) );
  CFA1X1 U438 ( .A(n467), .B(n490), .CI(n465), .CO(n460), .S(n461) );
  CFA1X1 U440 ( .A(n473), .B(n471), .CI(n496), .CO(n464), .S(n465) );
  CFA1X1 U441 ( .A(n475), .B(n498), .CI(n500), .CO(n466), .S(n467) );
  CFA1X1 U442 ( .A(n481), .B(n477), .CI(n479), .CO(n468), .S(n469) );
  CFA1X1 U443 ( .A(n502), .B(n483), .CI(n504), .CO(n470), .S(n471) );
  CFA1X1 U444 ( .A(n510), .B(n506), .CI(n508), .CO(n472), .S(n473) );
  CFA1X1 U445 ( .A(n1024), .B(n485), .CI(n1108), .CO(n474), .S(n475) );
  CFA1X1 U447 ( .A(n870), .B(n1078), .CI(n958), .CO(n478), .S(n479) );
  CFA1X1 U448 ( .A(n898), .B(n978), .CI(n924), .CO(n480), .S(n481) );
  CFA1X1 U449 ( .A(n880), .B(n910), .CI(n851), .CO(n482), .S(n483) );
  CHA1X1 U450 ( .A(n874), .B(n888), .CO(n484), .S(n485) );
  CFA1X1 U452 ( .A(n495), .B(n516), .CI(n493), .CO(n488), .S(n489) );
  CFA1X1 U453 ( .A(n497), .B(n518), .CI(n520), .CO(n490), .S(n491) );
  CFA1X1 U454 ( .A(n522), .B(n499), .CI(n501), .CO(n492), .S(n493) );
  CFA1X1 U455 ( .A(n503), .B(n524), .CI(n526), .CO(n494), .S(n495) );
  CFA1X1 U456 ( .A(n509), .B(n505), .CI(n507), .CO(n496), .S(n497) );
  CFA1X1 U457 ( .A(n530), .B(n511), .CI(n528), .CO(n498), .S(n499) );
  CFA1X1 U458 ( .A(n536), .B(n532), .CI(n534), .CO(n500), .S(n501) );
  CFA1X1 U459 ( .A(n979), .B(n1079), .CI(n1001), .CO(n502), .S(n503) );
  CFA1X1 U460 ( .A(n959), .B(n1051), .CI(n1109), .CO(n504), .S(n505) );
  CFA1X1 U461 ( .A(n911), .B(n1025), .CI(n925), .CO(n506), .S(n507) );
  CFA1X1 U462 ( .A(n889), .B(n941), .CI(n899), .CO(n508), .S(n509) );
  CFA1X1 U463 ( .A(n871), .B(n881), .CI(n875), .CO(n510), .S(n511) );
  CFA1X1 U464 ( .A(n517), .B(n515), .CI(n540), .CO(n512), .S(n513) );
  CFA1X1 U465 ( .A(n521), .B(n542), .CI(n519), .CO(n514), .S(n515) );
  CFA1X1 U466 ( .A(n546), .B(n544), .CI(n523), .CO(n516), .S(n517) );
  CFA1X1 U467 ( .A(n527), .B(n525), .CI(n548), .CO(n518), .S(n519) );
  CFA1X1 U468 ( .A(n533), .B(n550), .CI(n529), .CO(n520), .S(n521) );
  CFA1X1 U469 ( .A(n535), .B(n531), .CI(n552), .CO(n522), .S(n523) );
  CFA1X1 U470 ( .A(n558), .B(n554), .CI(n556), .CO(n524), .S(n525) );
  CFA1X1 U471 ( .A(n1002), .B(n560), .CI(n537), .CO(n526), .S(n527) );
  CFA1X1 U472 ( .A(n980), .B(n1080), .CI(n1110), .CO(n528), .S(n529) );
  CFA1X1 U473 ( .A(n926), .B(n1052), .CI(n960), .CO(n530), .S(n531) );
  CFA1X1 U474 ( .A(n912), .B(n1026), .CI(n876), .CO(n532), .S(n533) );
  CFA1X1 U475 ( .A(n890), .B(n900), .CI(n942), .CO(n534), .S(n535) );
  CHA1X1 U476 ( .A(n882), .B(n852), .CO(n536), .S(n537) );
  CFA1X1 U477 ( .A(n543), .B(n541), .CI(n564), .CO(n538), .S(n539) );
  CFA1X1 U478 ( .A(n568), .B(n566), .CI(n545), .CO(n540), .S(n541) );
  CFA1X1 U479 ( .A(n570), .B(n547), .CI(n549), .CO(n542), .S(n543) );
  CFA1X1 U480 ( .A(n574), .B(n551), .CI(n572), .CO(n544), .S(n545) );
  CFA1X1 U481 ( .A(n557), .B(n553), .CI(n555), .CO(n546), .S(n547) );
  CFA1X1 U482 ( .A(n578), .B(n559), .CI(n561), .CO(n548), .S(n549) );
  CFA1X1 U483 ( .A(n582), .B(n576), .CI(n580), .CO(n550), .S(n551) );
  CFA1X1 U484 ( .A(n1003), .B(n584), .CI(n1081), .CO(n552), .S(n553) );
  CFA1X1 U485 ( .A(n961), .B(n1053), .CI(n1111), .CO(n554), .S(n555) );
  CFA1X1 U486 ( .A(n913), .B(n1027), .CI(n1623), .CO(n556), .S(n557) );
  CFA1X1 U487 ( .A(n981), .B(n901), .CI(n927), .CO(n558), .S(n559) );
  CFA1X1 U488 ( .A(n877), .B(n891), .CI(n883), .CO(n560), .S(n561) );
  CFA1X1 U489 ( .A(n567), .B(n565), .CI(n588), .CO(n562), .S(n563) );
  CFA1X1 U490 ( .A(n592), .B(n590), .CI(n569), .CO(n564), .S(n565) );
  CFA1X1 U491 ( .A(n594), .B(n571), .CI(n573), .CO(n566), .S(n567) );
  CFA1X1 U492 ( .A(n598), .B(n575), .CI(n596), .CO(n568), .S(n569) );
  CFA1X1 U493 ( .A(n581), .B(n577), .CI(n579), .CO(n570), .S(n571) );
  CFA1X1 U494 ( .A(n602), .B(n583), .CI(n600), .CO(n572), .S(n573) );
  CFA1X1 U495 ( .A(n585), .B(n604), .CI(n606), .CO(n574), .S(n575) );
  CFA1X1 U496 ( .A(n1112), .B(n1004), .CI(n1028), .CO(n576), .S(n577) );
  CFA1X1 U497 ( .A(n884), .B(n1054), .CI(n982), .CO(n578), .S(n579) );
  CFA1X1 U498 ( .A(n928), .B(n1082), .CI(n962), .CO(n580), .S(n581) );
  CFA1X1 U499 ( .A(n853), .B(n1603), .CI(n914), .CO(n582), .S(n583) );
  CHA1X1 U500 ( .A(n892), .B(n902), .CO(n584), .S(n585) );
  CFA1X1 U502 ( .A(n614), .B(n612), .CI(n593), .CO(n588), .S(n589) );
  CFA1X1 U503 ( .A(n616), .B(n595), .CI(n597), .CO(n590), .S(n591) );
  CFA1X1 U504 ( .A(n601), .B(n599), .CI(n618), .CO(n592), .S(n593) );
  CFA1X1 U505 ( .A(n605), .B(n620), .CI(n603), .CO(n594), .S(n595) );
  CFA1X1 U506 ( .A(n624), .B(n607), .CI(n622), .CO(n596), .S(n597) );
  CFA1X1 U507 ( .A(n1005), .B(n626), .CI(n628), .CO(n598), .S(n599) );
  CFA1X1 U508 ( .A(n983), .B(n1055), .CI(n1113), .CO(n600), .S(n601) );
  CFA1X1 U509 ( .A(n929), .B(n1601), .CI(n963), .CO(n602), .S(n603) );
  CFA1X1 U510 ( .A(n915), .B(n1029), .CI(n1621), .CO(n604), .S(n605) );
  CFA1X1 U511 ( .A(n885), .B(n903), .CI(n893), .CO(n606), .S(n607) );
  CFA1X1 U512 ( .A(n613), .B(n611), .CI(n632), .CO(n608), .S(n609) );
  CFA1X1 U513 ( .A(n617), .B(n634), .CI(n615), .CO(n610), .S(n611) );
  CFA1X1 U514 ( .A(n638), .B(n636), .CI(n619), .CO(n612), .S(n613) );
  CFA1X1 U515 ( .A(n623), .B(n640), .CI(n621), .CO(n614), .S(n615) );
  CFA1X1 U516 ( .A(n642), .B(n625), .CI(n627), .CO(n616), .S(n617) );
  CFA1X1 U517 ( .A(n648), .B(n644), .CI(n646), .CO(n618), .S(n619) );
  CFA1X1 U518 ( .A(n1557), .B(n629), .CI(n1114), .CO(n620), .S(n621) );
  CFA1X1 U519 ( .A(n1616), .B(n1056), .CI(n1006), .CO(n622), .S(n623) );
  CFA1X1 U520 ( .A(n894), .B(n1084), .CI(n964), .CO(n624), .S(n625) );
  CFA1X1 U521 ( .A(n904), .B(n984), .CI(n930), .CO(n626), .S(n627) );
  CHA1X1 U522 ( .A(n854), .B(n916), .CO(n628), .S(n629) );
  CFA1X1 U523 ( .A(n635), .B(n633), .CI(n652), .CO(n630), .S(n631) );
  CFA1X1 U524 ( .A(n639), .B(n654), .CI(n637), .CO(n632), .S(n633) );
  CFA1X1 U525 ( .A(n658), .B(n656), .CI(n641), .CO(n634), .S(n635) );
  CFA1X1 U526 ( .A(n645), .B(n660), .CI(n643), .CO(n636), .S(n637) );
  CFA1X1 U527 ( .A(n662), .B(n647), .CI(n649), .CO(n638), .S(n639) );
  CFA1X1 U528 ( .A(n668), .B(n664), .CI(n666), .CO(n640), .S(n641) );
  CFA1X1 U530 ( .A(n1619), .B(n1085), .CI(n1007), .CO(n644), .S(n645) );
  CFA1X1 U531 ( .A(n931), .B(n1057), .CI(n965), .CO(n646), .S(n647) );
  CFA1X1 U532 ( .A(n895), .B(n917), .CI(n905), .CO(n648), .S(n649) );
  CFA1X1 U534 ( .A(n659), .B(n674), .CI(n657), .CO(n652), .S(n653) );
  CFA1X1 U535 ( .A(n678), .B(n676), .CI(n661), .CO(n654), .S(n655) );
  CFA1X1 U536 ( .A(n680), .B(n663), .CI(n665), .CO(n656), .S(n657) );
  CFA1X1 U537 ( .A(n684), .B(n667), .CI(n682), .CO(n658), .S(n659) );
  CFA1X1 U538 ( .A(n1008), .B(n686), .CI(n669), .CO(n660), .S(n661) );
  CFA1X1 U539 ( .A(n986), .B(n1086), .CI(n1116), .CO(n662), .S(n663) );
  CFA1X1 U540 ( .A(n932), .B(n966), .CI(n1058), .CO(n664), .S(n665) );
  CFA1X1 U541 ( .A(n918), .B(n1032), .CI(n948), .CO(n666), .S(n667) );
  CHA1X1 U542 ( .A(n855), .B(n906), .CO(n668), .S(n669) );
  CFA1X1 U543 ( .A(n675), .B(n673), .CI(n690), .CO(n670), .S(n671) );
  CFA1X1 U544 ( .A(n679), .B(n692), .CI(n677), .CO(n672), .S(n673) );
  CFA1X1 U545 ( .A(n681), .B(n694), .CI(n696), .CO(n674), .S(n675) );
  CFA1X1 U546 ( .A(n687), .B(n683), .CI(n685), .CO(n676), .S(n677) );
  CFA1X1 U547 ( .A(n702), .B(n698), .CI(n700), .CO(n678), .S(n679) );
  CFA1X1 U548 ( .A(n987), .B(n704), .CI(n1033), .CO(n680), .S(n681) );
  CFA1X1 U549 ( .A(n1087), .B(n967), .CI(n1117), .CO(n682), .S(n683) );
  CFA1X1 U550 ( .A(n949), .B(n1059), .CI(n1009), .CO(n684), .S(n685) );
  CFA1X1 U551 ( .A(n907), .B(n933), .CI(n919), .CO(n686), .S(n687) );
  CFA1X1 U552 ( .A(n693), .B(n691), .CI(n708), .CO(n688), .S(n689) );
  CFA1X1 U553 ( .A(n697), .B(n710), .CI(n695), .CO(n690), .S(n691) );
  CFA1X1 U554 ( .A(n699), .B(n712), .CI(n714), .CO(n692), .S(n693) );
  CFA1X1 U555 ( .A(n718), .B(n701), .CI(n703), .CO(n694), .S(n695) );
  CFA1X1 U556 ( .A(n705), .B(n716), .CI(n720), .CO(n696), .S(n697) );
  CFA1X1 U557 ( .A(n1010), .B(n1118), .CI(n1034), .CO(n698), .S(n699) );
  CFA1X1 U558 ( .A(n920), .B(n1088), .CI(n988), .CO(n700), .S(n701) );
  CFA1X1 U559 ( .A(n934), .B(n968), .CI(n1612), .CO(n702), .S(n703) );
  CHA1X1 U560 ( .A(n856), .B(n950), .CO(n704), .S(n705) );
  CFA1X1 U561 ( .A(n711), .B(n709), .CI(n724), .CO(n706), .S(n707) );
  CFA1X1 U562 ( .A(n715), .B(n726), .CI(n713), .CO(n708), .S(n709) );
  CFA1X1 U563 ( .A(n717), .B(n728), .CI(n730), .CO(n710), .S(n711) );
  CFA1X1 U564 ( .A(n732), .B(n719), .CI(n721), .CO(n712), .S(n713) );
  CFA1X1 U565 ( .A(n1011), .B(n734), .CI(n736), .CO(n714), .S(n715) );
  CFA1X1 U566 ( .A(n989), .B(n1089), .CI(n1035), .CO(n716), .S(n717) );
  CFA1X1 U567 ( .A(n969), .B(n1061), .CI(n1119), .CO(n718), .S(n719) );
  CFA1X1 U568 ( .A(n921), .B(n951), .CI(n935), .CO(n720), .S(n721) );
  CFA1X1 U569 ( .A(n727), .B(n725), .CI(n740), .CO(n722), .S(n723) );
  CFA1X1 U570 ( .A(n744), .B(n742), .CI(n729), .CO(n724), .S(n725) );
  CFA1X1 U571 ( .A(n735), .B(n731), .CI(n733), .CO(n726), .S(n727) );
  CFA1X1 U572 ( .A(n750), .B(n748), .CI(n746), .CO(n728), .S(n729) );
  CFA1X1 U573 ( .A(n970), .B(n737), .CI(n1120), .CO(n730), .S(n731) );
  CFA1X1 U574 ( .A(n1561), .B(n1090), .CI(n1036), .CO(n732), .S(n733) );
  CFA1X1 U575 ( .A(n1625), .B(n1062), .CI(n1012), .CO(n734), .S(n735) );
  CFA1X1 U577 ( .A(n743), .B(n741), .CI(n754), .CO(n738), .S(n739) );
  CFA1X1 U578 ( .A(n758), .B(n756), .CI(n745), .CO(n740), .S(n741) );
  CFA1X1 U579 ( .A(n751), .B(n747), .CI(n749), .CO(n742), .S(n743) );
  CFA1X1 U580 ( .A(n764), .B(n762), .CI(n760), .CO(n744), .S(n745) );
  CFA1X1 U581 ( .A(n1013), .B(n1121), .CI(n1037), .CO(n746), .S(n747) );
  CFA1X1 U582 ( .A(n991), .B(n1091), .CI(n1063), .CO(n748), .S(n749) );
  CFA1X1 U583 ( .A(n937), .B(n971), .CI(n953), .CO(n750), .S(n751) );
  CFA1X1 U584 ( .A(n757), .B(n755), .CI(n768), .CO(n752), .S(n753) );
  CFA1X1 U585 ( .A(n772), .B(n759), .CI(n770), .CO(n754), .S(n755) );
  CFA1X1 U586 ( .A(n774), .B(n761), .CI(n763), .CO(n756), .S(n757) );
  CFA1X1 U587 ( .A(n992), .B(n776), .CI(n765), .CO(n758), .S(n759) );
  CFA1X1 U589 ( .A(n972), .B(n1064), .CI(n1122), .CO(n762), .S(n763) );
  CHA1X1 U590 ( .A(n858), .B(n1014), .CO(n764), .S(n765) );
  CFA1X1 U591 ( .A(n771), .B(n769), .CI(n780), .CO(n766), .S(n767) );
  CFA1X1 U592 ( .A(n775), .B(n782), .CI(n773), .CO(n768), .S(n769) );
  CFA1X1 U593 ( .A(n784), .B(n777), .CI(n786), .CO(n770), .S(n771) );
  CFA1X1 U595 ( .A(n1558), .B(n1065), .CI(n1093), .CO(n774), .S(n775) );
  CFA1X1 U596 ( .A(n955), .B(n993), .CI(n973), .CO(n776), .S(n777) );
  CFA1X1 U597 ( .A(n783), .B(n781), .CI(n792), .CO(n778), .S(n779) );
  CFA1X1 U598 ( .A(n787), .B(n794), .CI(n785), .CO(n780), .S(n781) );
  CFA1X1 U599 ( .A(n789), .B(n796), .CI(n798), .CO(n782), .S(n783) );
  CFA1X1 U600 ( .A(n994), .B(n1040), .CI(n1016), .CO(n784), .S(n785) );
  CFA1X1 U601 ( .A(n974), .B(n1066), .CI(n1124), .CO(n786), .S(n787) );
  CFA1X1 U603 ( .A(n802), .B(n793), .CI(n795), .CO(n790), .S(n791) );
  CFA1X1 U604 ( .A(n799), .B(n804), .CI(n797), .CO(n792), .S(n793) );
  CFA1X1 U605 ( .A(n1125), .B(n806), .CI(n808), .CO(n794), .S(n795) );
  CFA1X1 U607 ( .A(n975), .B(n1017), .CI(n1559), .CO(n798), .S(n799) );
  CFA1X1 U608 ( .A(n805), .B(n803), .CI(n812), .CO(n800), .S(n801) );
  CFA1X1 U609 ( .A(n816), .B(n807), .CI(n814), .CO(n802), .S(n803) );
  CFA1X1 U610 ( .A(n1018), .B(n809), .CI(n1042), .CO(n804), .S(n805) );
  CFA1X1 U611 ( .A(n996), .B(n1068), .CI(n1126), .CO(n806), .S(n807) );
  CHA1X1 U612 ( .A(n860), .B(n1096), .CO(n808), .S(n809) );
  CFA1X1 U613 ( .A(n815), .B(n813), .CI(n820), .CO(n810), .S(n811) );
  CFA1X1 U614 ( .A(n824), .B(n817), .CI(n822), .CO(n812), .S(n813) );
  CFA1X1 U615 ( .A(n1127), .B(n1097), .CI(n1069), .CO(n814), .S(n815) );
  CFA1X1 U617 ( .A(n828), .B(n821), .CI(n823), .CO(n818), .S(n819) );
  CFA1X1 U618 ( .A(n1044), .B(n830), .CI(n825), .CO(n820), .S(n821) );
  CFA1X1 U619 ( .A(n1020), .B(n1070), .CI(n1128), .CO(n822), .S(n823) );
  CHA1X1 U620 ( .A(n861), .B(n1098), .CO(n824), .S(n825) );
  CFA1X1 U621 ( .A(n834), .B(n829), .CI(n831), .CO(n826), .S(n827) );
  CFA1X1 U622 ( .A(n1099), .B(n836), .CI(n1071), .CO(n828), .S(n829) );
  CFA1X1 U624 ( .A(n837), .B(n835), .CI(n840), .CO(n832), .S(n833) );
  CFA1X1 U625 ( .A(n1046), .B(n1072), .CI(n1130), .CO(n834), .S(n835) );
  CHA1X1 U626 ( .A(n862), .B(n1100), .CO(n836), .S(n837) );
  CFA1X1 U627 ( .A(n1073), .B(n841), .CI(n844), .CO(n838), .S(n839) );
  CFA1X1 U628 ( .A(n1047), .B(n1101), .CI(n1131), .CO(n840), .S(n841) );
  CFA1X1 U629 ( .A(n1102), .B(n845), .CI(n1074), .CO(n842), .S(n843) );
  CHA1X1 U630 ( .A(n1132), .B(n863), .CO(n844), .S(n845) );
  CFA1X1 U631 ( .A(n1075), .B(n1103), .CI(n1133), .CO(n846), .S(n847) );
  CHA1X1 U632 ( .A(n1134), .B(n1104), .CO(n848), .S(n849) );
  COND2X1 U633 ( .A(n115), .B(n1468), .C(n114), .D(n1139), .Z(n850) );
  COND2X1 U634 ( .A(n1138), .B(n115), .C(n114), .D(n1137), .Z(n866) );
  CND2IX1 U638 ( .B(n1746), .A(n113), .Z(n1139) );
  COND2X1 U639 ( .A(n112), .B(n1469), .C(n110), .D(n1144), .Z(n851) );
  COND2X1 U640 ( .A(n112), .B(n1141), .C(n110), .D(n1140), .Z(n868) );
  COND2X1 U642 ( .A(n1143), .B(n112), .C(n110), .D(n1142), .Z(n870) );
  CND2IX1 U648 ( .B(n1746), .A(n109), .Z(n1144) );
  COND2X1 U649 ( .A(n1151), .B(n105), .C(n1470), .D(n107), .Z(n852) );
  COND2X1 U651 ( .A(n107), .B(n1147), .C(n105), .D(n1146), .Z(n873) );
  COND2X1 U653 ( .A(n107), .B(n1149), .C(n105), .D(n1148), .Z(n875) );
  COND2X1 U654 ( .A(n1150), .B(n107), .C(n105), .D(n1149), .Z(n876) );
  CND2IX1 U662 ( .B(n1746), .A(n1717), .Z(n1151) );
  COND2X1 U663 ( .A(n102), .B(n1591), .C(n100), .D(n1160), .Z(n853) );
  COND2X1 U664 ( .A(n102), .B(n1153), .C(n100), .D(n1152), .Z(n878) );
  COND2X1 U665 ( .A(n102), .B(n1154), .C(n100), .D(n1153), .Z(n879) );
  COND2X1 U666 ( .A(n102), .B(n1155), .C(n100), .D(n1154), .Z(n880) );
  COND2X1 U667 ( .A(n102), .B(n1156), .C(n100), .D(n1155), .Z(n881) );
  COND2X1 U668 ( .A(n102), .B(n1157), .C(n100), .D(n1156), .Z(n882) );
  COND2X1 U669 ( .A(n102), .B(n1158), .C(n100), .D(n1157), .Z(n883) );
  COND2X1 U670 ( .A(n1159), .B(n102), .C(n100), .D(n1158), .Z(n884) );
  CND2IX1 U680 ( .B(n1746), .A(n1716), .Z(n1160) );
  COND2X1 U681 ( .A(n97), .B(n1472), .C(n95), .D(n1171), .Z(n854) );
  COND2X1 U686 ( .A(n97), .B(n1166), .C(n1165), .D(n95), .Z(n890) );
  COND2X1 U687 ( .A(n97), .B(n1167), .C(n1166), .D(n95), .Z(n891) );
  COND2X1 U703 ( .A(n91), .B(n1473), .C(n1563), .D(n1184), .Z(n855) );
  COND2X1 U704 ( .A(n91), .B(n1173), .C(n1172), .D(n1563), .Z(n896) );
  COND2X1 U705 ( .A(n91), .B(n1174), .C(n1173), .D(n1563), .Z(n897) );
  COND2X1 U706 ( .A(n91), .B(n1175), .C(n1174), .D(n1563), .Z(n898) );
  COND2X1 U707 ( .A(n91), .B(n1176), .C(n1175), .D(n1604), .Z(n899) );
  COND2X1 U708 ( .A(n91), .B(n1177), .C(n1176), .D(n1563), .Z(n900) );
  COND2X1 U709 ( .A(n91), .B(n1178), .C(n1177), .D(n1604), .Z(n901) );
  COND2X1 U710 ( .A(n91), .B(n1179), .C(n1178), .D(n1604), .Z(n902) );
  COND2X1 U711 ( .A(n91), .B(n1180), .C(n1179), .D(n1604), .Z(n903) );
  COND2X1 U712 ( .A(n91), .B(n1181), .C(n1180), .D(n1563), .Z(n904) );
  COND2X1 U713 ( .A(n91), .B(n1182), .C(n1181), .D(n1604), .Z(n905) );
  COND2X1 U714 ( .A(n1183), .B(n91), .C(n1182), .D(n1604), .Z(n906) );
  CND2IX1 U728 ( .B(n1746), .A(n1714), .Z(n1184) );
  COND2X1 U732 ( .A(n85), .B(n1188), .C(n1187), .D(n82), .Z(n910) );
  COND2X1 U734 ( .A(n85), .B(n1190), .C(n1189), .D(n82), .Z(n912) );
  COND2X1 U735 ( .A(n85), .B(n1191), .C(n1190), .D(n82), .Z(n913) );
  COND2X1 U736 ( .A(n85), .B(n1192), .C(n1191), .D(n82), .Z(n914) );
  COND2X1 U737 ( .A(n85), .B(n1193), .C(n1192), .D(n82), .Z(n915) );
  COND2X1 U739 ( .A(n85), .B(n1195), .C(n1194), .D(n82), .Z(n917) );
  COND2X1 U740 ( .A(n85), .B(n1196), .C(n1195), .D(n82), .Z(n918) );
  COND2X1 U741 ( .A(n85), .B(n1197), .C(n1196), .D(n82), .Z(n919) );
  CND2IX1 U758 ( .B(n1746), .A(n1713), .Z(n1199) );
  COND2X1 U761 ( .A(n77), .B(n1202), .C(n1201), .D(n74), .Z(n923) );
  COND2X1 U762 ( .A(n77), .B(n1203), .C(n1202), .D(n74), .Z(n924) );
  COND2X1 U763 ( .A(n77), .B(n1204), .C(n1203), .D(n74), .Z(n925) );
  COND2X1 U765 ( .A(n77), .B(n1206), .C(n1205), .D(n74), .Z(n927) );
  COND2X1 U766 ( .A(n77), .B(n1207), .C(n1206), .D(n74), .Z(n928) );
  COND2X1 U767 ( .A(n77), .B(n1208), .C(n1207), .D(n74), .Z(n929) );
  COND2X1 U768 ( .A(n77), .B(n1209), .C(n1208), .D(n74), .Z(n930) );
  COND2X1 U769 ( .A(n77), .B(n1210), .C(n1209), .D(n74), .Z(n931) );
  COND2X1 U770 ( .A(n77), .B(n1211), .C(n1210), .D(n74), .Z(n932) );
  COND2X1 U771 ( .A(n77), .B(n1212), .C(n1211), .D(n74), .Z(n933) );
  COND2X1 U773 ( .A(n77), .B(n1214), .C(n1213), .D(n74), .Z(n935) );
  COND2X1 U798 ( .A(n69), .B(n1222), .C(n1221), .D(n66), .Z(n942) );
  COND2X1 U804 ( .A(n69), .B(n1228), .C(n1227), .D(n66), .Z(n948) );
  COND2X1 U805 ( .A(n69), .B(n1229), .C(n1228), .D(n66), .Z(n949) );
  COND2X1 U806 ( .A(n69), .B(n1230), .C(n1229), .D(n66), .Z(n950) );
  COND2X1 U807 ( .A(n69), .B(n1231), .C(n1230), .D(n66), .Z(n951) );
  COND2X1 U809 ( .A(n69), .B(n1233), .C(n1232), .D(n66), .Z(n953) );
  COND2X1 U832 ( .A(n61), .B(n1237), .C(n1236), .D(n1617), .Z(n956) );
  COND2X1 U833 ( .A(n61), .B(n1238), .C(n1237), .D(n1617), .Z(n957) );
  COND2X1 U834 ( .A(n61), .B(n1239), .C(n1238), .D(n1617), .Z(n958) );
  COND2X1 U835 ( .A(n61), .B(n1240), .C(n1239), .D(n1617), .Z(n959) );
  COND2X1 U836 ( .A(n61), .B(n1241), .C(n1240), .D(n1617), .Z(n960) );
  COND2X1 U837 ( .A(n61), .B(n1242), .C(n1241), .D(n1617), .Z(n961) );
  COND2X1 U838 ( .A(n61), .B(n1243), .C(n1242), .D(n1617), .Z(n962) );
  COND2X1 U839 ( .A(n61), .B(n1244), .C(n1243), .D(n1617), .Z(n963) );
  COND2X1 U840 ( .A(n61), .B(n1245), .C(n1244), .D(n1617), .Z(n964) );
  COND2X1 U841 ( .A(n61), .B(n1246), .C(n1245), .D(n1617), .Z(n965) );
  COND2X1 U842 ( .A(n61), .B(n1247), .C(n1246), .D(n1617), .Z(n966) );
  COND2X1 U843 ( .A(n61), .B(n1248), .C(n1247), .D(n1617), .Z(n967) );
  COND2X1 U844 ( .A(n61), .B(n1249), .C(n1248), .D(n1617), .Z(n968) );
  COND2X1 U845 ( .A(n61), .B(n1250), .C(n1249), .D(n1617), .Z(n969) );
  COND2X1 U846 ( .A(n61), .B(n1251), .C(n1250), .D(n1617), .Z(n970) );
  COND2X1 U847 ( .A(n61), .B(n1252), .C(n1251), .D(n1617), .Z(n971) );
  COND2X1 U848 ( .A(n61), .B(n1253), .C(n1252), .D(n1617), .Z(n972) );
  COND2X1 U849 ( .A(n61), .B(n1254), .C(n1253), .D(n1617), .Z(n973) );
  COND2X1 U850 ( .A(n61), .B(n1255), .C(n1254), .D(n1617), .Z(n974) );
  COND2X1 U878 ( .A(n53), .B(n1262), .C(n1261), .D(n50), .Z(n980) );
  COND2X1 U879 ( .A(n53), .B(n1263), .C(n1262), .D(n50), .Z(n981) );
  COND2X1 U884 ( .A(n53), .B(n1268), .C(n1267), .D(n50), .Z(n986) );
  COND2X1 U886 ( .A(n53), .B(n1270), .C(n1269), .D(n50), .Z(n988) );
  COND2X1 U889 ( .A(n53), .B(n1273), .C(n1272), .D(n50), .Z(n991) );
  COND2X1 U923 ( .A(n44), .B(n1284), .C(n1283), .D(n1654), .Z(n1001) );
  COND2X1 U925 ( .A(n44), .B(n1286), .C(n1285), .D(n1654), .Z(n1003) );
  COND2X1 U928 ( .A(n44), .B(n1289), .C(n1288), .D(n1654), .Z(n1006) );
  COND2X1 U929 ( .A(n44), .B(n1290), .C(n1289), .D(n1654), .Z(n1007) );
  COND2X1 U931 ( .A(n44), .B(n1292), .C(n1291), .D(n1654), .Z(n1009) );
  COND2X1 U932 ( .A(n44), .B(n1293), .C(n1292), .D(n1654), .Z(n1010) );
  COND2X1 U934 ( .A(n44), .B(n1295), .C(n1294), .D(n1654), .Z(n1012) );
  COND2X1 U935 ( .A(n44), .B(n1296), .C(n1295), .D(n1654), .Z(n1013) );
  COND2X1 U936 ( .A(n44), .B(n1297), .C(n1296), .D(n1654), .Z(n1014) );
  COND2X1 U938 ( .A(n44), .B(n1299), .C(n1298), .D(n1654), .Z(n1016) );
  COND2X1 U939 ( .A(n44), .B(n1300), .C(n1299), .D(n1654), .Z(n1017) );
  COND2X1 U941 ( .A(n44), .B(n1302), .C(n1301), .D(n1654), .Z(n1019) );
  CND2IX1 U968 ( .B(n1746), .A(n1740), .Z(n1304) );
  COND2X1 U975 ( .A(n36), .B(n1311), .C(n1310), .D(n1658), .Z(n1027) );
  COND2X1 U980 ( .A(n36), .B(n1316), .C(n1315), .D(n1658), .Z(n1032) );
  COND2X1 U982 ( .A(n36), .B(n1318), .C(n1317), .D(n1658), .Z(n1034) );
  COND2X1 U984 ( .A(n36), .B(n1320), .C(n1319), .D(n1658), .Z(n1036) );
  COND2X1 U985 ( .A(n36), .B(n1321), .C(n1320), .D(n1658), .Z(n1037) );
  COND2X1 U986 ( .A(n36), .B(n1322), .C(n1321), .D(n1658), .Z(n1038) );
  COND2X1 U1028 ( .A(n27), .B(n1337), .C(n1653), .D(n1336), .Z(n1052) );
  COND2X1 U1035 ( .A(n27), .B(n1344), .C(n1653), .D(n1343), .Z(n1059) );
  COND2X1 U1037 ( .A(n27), .B(n1346), .C(n1653), .D(n1345), .Z(n1061) );
  COND2X1 U1039 ( .A(n27), .B(n1348), .C(n1653), .D(n1347), .Z(n1063) );
  COND2X1 U1040 ( .A(n27), .B(n1349), .C(n1653), .D(n1348), .Z(n1064) );
  COND2X1 U1043 ( .A(n27), .B(n1352), .C(n1653), .D(n1351), .Z(n1067) );
  CND2IX1 U1080 ( .B(n1746), .A(n1727), .Z(n1360) );
  COND2X1 U1086 ( .A(n18), .B(n1366), .C(n1631), .D(n1365), .Z(n1080) );
  COND2X1 U1087 ( .A(n18), .B(n1367), .C(n1632), .D(n1366), .Z(n1081) );
  COND2X1 U1088 ( .A(n18), .B(n1368), .C(n1631), .D(n1367), .Z(n1082) );
  COND2X1 U1091 ( .A(n18), .B(n1371), .C(n1632), .D(n1370), .Z(n1085) );
  COND2X1 U1092 ( .A(n18), .B(n1372), .C(n1632), .D(n1371), .Z(n1086) );
  COND2X1 U1094 ( .A(n18), .B(n1374), .C(n1631), .D(n1373), .Z(n1088) );
  COND2X1 U1096 ( .A(n18), .B(n1376), .C(n1631), .D(n1375), .Z(n1090) );
  COND2X1 U1097 ( .A(n18), .B(n1377), .C(n1632), .D(n1376), .Z(n1091) );
  COND2X1 U1098 ( .A(n18), .B(n1378), .C(n1632), .D(n1377), .Z(n1092) );
  COND2X1 U1100 ( .A(n18), .B(n1380), .C(n1632), .D(n1379), .Z(n1094) );
  COND2X1 U1102 ( .A(n18), .B(n1382), .C(n1631), .D(n1381), .Z(n1096) );
  CND2IX1 U1142 ( .B(n1746), .A(n1719), .Z(n1391) );
  COND2X1 U1144 ( .A(n9), .B(n1393), .C(n6), .D(n1392), .Z(n1106) );
  COND2X1 U1145 ( .A(n9), .B(n1394), .C(n6), .D(n1393), .Z(n1107) );
  COND2X1 U1146 ( .A(n9), .B(n1395), .C(n6), .D(n1394), .Z(n1108) );
  COND2X1 U1147 ( .A(n9), .B(n1396), .C(n6), .D(n1395), .Z(n1109) );
  COND2X1 U1148 ( .A(n9), .B(n1397), .C(n6), .D(n1396), .Z(n1110) );
  COND2X1 U1149 ( .A(n9), .B(n1398), .C(n6), .D(n1397), .Z(n1111) );
  COND2X1 U1150 ( .A(n9), .B(n1399), .C(n6), .D(n1398), .Z(n1112) );
  COND2X1 U1151 ( .A(n9), .B(n1400), .C(n6), .D(n1399), .Z(n1113) );
  COND2X1 U1152 ( .A(n9), .B(n1401), .C(n6), .D(n1400), .Z(n1114) );
  COND2X1 U1153 ( .A(n9), .B(n1402), .C(n6), .D(n1401), .Z(n1115) );
  COND2X1 U1154 ( .A(n9), .B(n1403), .C(n6), .D(n1402), .Z(n1116) );
  COND2X1 U1155 ( .A(n9), .B(n1404), .C(n6), .D(n1403), .Z(n1117) );
  COND2X1 U1156 ( .A(n9), .B(n1405), .C(n6), .D(n1404), .Z(n1118) );
  COND2X1 U1157 ( .A(n9), .B(n1406), .C(n6), .D(n1405), .Z(n1119) );
  COND2X1 U1158 ( .A(n9), .B(n1407), .C(n6), .D(n1406), .Z(n1120) );
  COND2X1 U1159 ( .A(n9), .B(n1408), .C(n6), .D(n1407), .Z(n1121) );
  COND2X1 U1160 ( .A(n9), .B(n1409), .C(n6), .D(n1408), .Z(n1122) );
  COND2X1 U1161 ( .A(n9), .B(n1410), .C(n6), .D(n1409), .Z(n1123) );
  COND2X1 U1162 ( .A(n9), .B(n1411), .C(n6), .D(n1410), .Z(n1124) );
  COND2X1 U1163 ( .A(n9), .B(n1412), .C(n6), .D(n1411), .Z(n1125) );
  COND2X1 U1164 ( .A(n9), .B(n1413), .C(n6), .D(n1412), .Z(n1126) );
  COND2X1 U1165 ( .A(n9), .B(n1414), .C(n6), .D(n1413), .Z(n1127) );
  COND2X1 U1166 ( .A(n9), .B(n1415), .C(n6), .D(n1414), .Z(n1128) );
  COND2X1 U1167 ( .A(n9), .B(n1416), .C(n6), .D(n1415), .Z(n1129) );
  COND2X1 U1168 ( .A(n9), .B(n1417), .C(n6), .D(n1416), .Z(n1130) );
  COND2X1 U1169 ( .A(n9), .B(n1418), .C(n6), .D(n1417), .Z(n1131) );
  COND2X1 U1170 ( .A(n9), .B(n1419), .C(n6), .D(n1418), .Z(n1132) );
  COND2X1 U1171 ( .A(n9), .B(n1420), .C(n6), .D(n1419), .Z(n1133) );
  COND2X1 U1172 ( .A(n9), .B(n1421), .C(n6), .D(n1420), .Z(n1134) );
  COND2X1 U1173 ( .A(n9), .B(n1422), .C(n6), .D(n1421), .Z(n1135) );
  COND2X1 U1174 ( .A(n9), .B(n1423), .C(n6), .D(n1422), .Z(n1136) );
  CND2IX1 U1208 ( .B(n1746), .A(n1718), .Z(n1424) );
  CENX1 U1281 ( .A(n1743), .B(n1701), .Z(n1272) );
  CENX1 U1282 ( .A(n1711), .B(n1701), .Z(n1228) );
  CENX1 U1283 ( .A(n1711), .B(n1697), .Z(n1232) );
  CENX1 U1284 ( .A(n1697), .B(n1717), .Z(n1148) );
  CANR1X2 U1285 ( .A(n229), .B(n216), .C(n217), .Z(n1575) );
  COND2X1 U1286 ( .A(n85), .B(n1187), .C(n1186), .D(n82), .Z(n909) );
  CIVX2 U1287 ( .A(n1060), .Z(n1611) );
  CENX1 U1288 ( .A(n1743), .B(n1696), .Z(n1277) );
  CENXL U1289 ( .A(n1712), .B(n1696), .Z(n1214) );
  CENXL U1290 ( .A(n1738), .B(n1696), .Z(n1302) );
  COND2X1 U1291 ( .A(n85), .B(n1474), .C(n82), .D(n1199), .Z(n856) );
  CND2X2 U1292 ( .A(n1666), .B(n1664), .Z(n245) );
  COND1X1 U1293 ( .A(n328), .B(n322), .C(n323), .Z(n321) );
  CNIVX1 U1294 ( .A(n1030), .Z(n1557) );
  CENXL U1295 ( .A(n1696), .B(n1717), .Z(n1149) );
  CNIVX3 U1296 ( .A(n104), .Z(n1717) );
  CNIVX1 U1297 ( .A(n1015), .Z(n1558) );
  CNIVX1 U1298 ( .A(n995), .Z(n1559) );
  CENXL U1299 ( .A(n1661), .B(n1703), .Z(n1415) );
  CENXL U1300 ( .A(n1723), .B(n1703), .Z(n1382) );
  CENXL U1301 ( .A(n1713), .B(n1703), .Z(n1190) );
  CENXL U1302 ( .A(n1682), .B(n1703), .Z(n1351) );
  CENX1 U1303 ( .A(n1743), .B(n1703), .Z(n1270) );
  COND2XL U1304 ( .A(n36), .B(n1314), .C(n1313), .D(n1658), .Z(n1030) );
  COND2XL U1305 ( .A(n36), .B(n1310), .C(n1309), .D(n1658), .Z(n1026) );
  COND2XL U1306 ( .A(n36), .B(n1317), .C(n1316), .D(n1658), .Z(n1033) );
  CENX1 U1307 ( .A(a[10]), .B(n1568), .Z(n1656) );
  CIVDX2 U1308 ( .A(n48), .Z0(n1567), .Z1(n1568) );
  CIVDX3 U1309 ( .A(n55), .Z0(n1569), .Z1(n1570) );
  CNIVX4 U1310 ( .A(n58), .Z(n1617) );
  CENXL U1311 ( .A(n1661), .B(n1705), .Z(n1413) );
  CENXL U1312 ( .A(n1739), .B(n1705), .Z(n1293) );
  CENXL U1313 ( .A(n1570), .B(n1705), .Z(n1245) );
  CENXL U1314 ( .A(n1682), .B(n1705), .Z(n1349) );
  CENXL U1315 ( .A(n1734), .B(n1705), .Z(n1320) );
  CENXL U1316 ( .A(n1713), .B(n1705), .Z(n1188) );
  CND2X4 U1317 ( .A(n1637), .B(n1638), .Z(n1653) );
  CND2X2 U1318 ( .A(n1635), .B(n1636), .Z(n1638) );
  CENXL U1319 ( .A(n1627), .B(n153), .Z(n1236) );
  CENXL U1320 ( .A(n1726), .B(n153), .Z(n1340) );
  CENXL U1321 ( .A(n1711), .B(n151), .Z(n1217) );
  CENXL U1322 ( .A(n1746), .B(n1711), .Z(n1234) );
  CENXL U1323 ( .A(n1711), .B(n1709), .Z(n1220) );
  CENXL U1324 ( .A(n1711), .B(n1703), .Z(n1226) );
  CENXL U1325 ( .A(n1711), .B(n1710), .Z(n1219) );
  CENXL U1326 ( .A(n1711), .B(n1708), .Z(n1221) );
  CENXL U1327 ( .A(n1711), .B(n1704), .Z(n1225) );
  CENXL U1328 ( .A(n1711), .B(n1699), .Z(n1230) );
  CENXL U1329 ( .A(n1711), .B(n1702), .Z(n1227) );
  CENXL U1330 ( .A(n1711), .B(n1700), .Z(n1229) );
  CENXL U1331 ( .A(n1711), .B(n1705), .Z(n1224) );
  CENXL U1332 ( .A(n1711), .B(n1698), .Z(n1231) );
  CENXL U1333 ( .A(n1711), .B(n1706), .Z(n1223) );
  CENXL U1334 ( .A(n1711), .B(n1707), .Z(n1222) );
  CND2XL U1335 ( .A(n1597), .B(n1711), .Z(n1599) );
  CENXL U1336 ( .A(n1743), .B(n155), .Z(n1257) );
  CENXL U1337 ( .A(n1743), .B(n1699), .Z(n1274) );
  CENXL U1338 ( .A(n1743), .B(n154), .Z(n1258) );
  CENXL U1339 ( .A(n1743), .B(n1700), .Z(n1273) );
  CENXL U1340 ( .A(n1743), .B(n1708), .Z(n1265) );
  CENXL U1341 ( .A(n1743), .B(n1698), .Z(n1275) );
  CENXL U1342 ( .A(n1743), .B(n1702), .Z(n1271) );
  CENXL U1343 ( .A(n1743), .B(n1697), .Z(n1276) );
  CIVX1 U1344 ( .A(n936), .Z(n1560) );
  CIVX2 U1345 ( .A(n1560), .Z(n1561) );
  CANR1X1 U1346 ( .A(n1677), .B(n357), .C(n354), .Z(n352) );
  COND1X1 U1347 ( .A(n358), .B(n360), .C(n359), .Z(n357) );
  COR2XL U1348 ( .A(n53), .B(n1264), .Z(n1587) );
  CNIVX1 U1349 ( .A(n1744), .Z(n1628) );
  CNIVX2 U1350 ( .A(n126), .Z(n1699) );
  CNIVX2 U1351 ( .A(n122), .Z(n1697) );
  CNIVX1 U1352 ( .A(n1744), .Z(n1627) );
  CNIVX1 U1353 ( .A(n148), .Z(n1710) );
  CND2X1 U1354 ( .A(n1598), .B(n1599), .Z(n1451) );
  CNIVX1 U1355 ( .A(n1744), .Z(n1626) );
  CENX1 U1356 ( .A(n1712), .B(n1698), .Z(n1212) );
  CENX1 U1357 ( .A(n1712), .B(n1697), .Z(n1213) );
  CENX1 U1358 ( .A(n1713), .B(n1696), .Z(n1197) );
  CENX1 U1359 ( .A(n1570), .B(n1702), .Z(n1248) );
  CENX1 U1360 ( .A(n1719), .B(n153), .Z(n1371) );
  CENX1 U1361 ( .A(n1570), .B(n1703), .Z(n1247) );
  CENX1 U1362 ( .A(n1712), .B(n1700), .Z(n1210) );
  CENX1 U1363 ( .A(n1712), .B(n1699), .Z(n1211) );
  CENX1 U1364 ( .A(n1712), .B(n1701), .Z(n1209) );
  CENX1 U1365 ( .A(n1730), .B(n152), .Z(n1341) );
  CENX1 U1366 ( .A(n1712), .B(n1702), .Z(n1208) );
  CENX1 U1367 ( .A(n1736), .B(n152), .Z(n1312) );
  CENX1 U1368 ( .A(n1570), .B(n1707), .Z(n1243) );
  CENX1 U1369 ( .A(n1712), .B(n1703), .Z(n1207) );
  CENX1 U1370 ( .A(n1712), .B(n1704), .Z(n1206) );
  CENX1 U1371 ( .A(n1723), .B(n1705), .Z(n1380) );
  CENX1 U1372 ( .A(n1570), .B(n1696), .Z(n1254) );
  CENX1 U1373 ( .A(n1723), .B(n1704), .Z(n1381) );
  CENX1 U1374 ( .A(n1570), .B(n1697), .Z(n1253) );
  CENX1 U1375 ( .A(n1746), .B(n1712), .Z(n1215) );
  CENX1 U1376 ( .A(n1570), .B(n1700), .Z(n1250) );
  CENX1 U1377 ( .A(n1724), .B(n150), .Z(n1374) );
  CND2X1 U1378 ( .A(n1587), .B(n1588), .Z(n982) );
  CNIVX2 U1379 ( .A(n130), .Z(n1701) );
  CNIVX1 U1380 ( .A(n138), .Z(n1705) );
  CND2X1 U1381 ( .A(a[14]), .B(n1639), .Z(n1598) );
  CENX1 U1382 ( .A(n1740), .B(n153), .Z(n1284) );
  CENX1 U1383 ( .A(n1712), .B(n1707), .Z(n1203) );
  CENX1 U1384 ( .A(n1696), .B(n109), .Z(n1142) );
  CND2X1 U1385 ( .A(n1581), .B(n1582), .Z(n926) );
  CENX1 U1386 ( .A(n1738), .B(n1698), .Z(n1300) );
  CENX1 U1387 ( .A(n1738), .B(n1697), .Z(n1301) );
  CNR2IX1 U1388 ( .B(n1746), .A(n74), .Z(n937) );
  CNIVX1 U1389 ( .A(n134), .Z(n1703) );
  CNIVX2 U1390 ( .A(n128), .Z(n1700) );
  CENX1 U1391 ( .A(n1743), .B(n153), .Z(n1259) );
  CENX1 U1392 ( .A(n1712), .B(n1708), .Z(n1202) );
  CNIVX2 U1393 ( .A(n99), .Z(n1716) );
  CNIVX4 U1394 ( .A(n79), .Z(n1713) );
  CND2X1 U1395 ( .A(n1644), .B(n1645), .Z(n1647) );
  CNIVX2 U1396 ( .A(n124), .Z(n1698) );
  CENX1 U1397 ( .A(n1697), .B(n109), .Z(n1141) );
  CND2IX2 U1398 ( .B(n1652), .A(n1653), .Z(n27) );
  CND2X1 U1399 ( .A(n1720), .B(a[4]), .Z(n1637) );
  CNIVX2 U1400 ( .A(n120), .Z(n1696) );
  CND2X2 U1401 ( .A(n1457), .B(n15), .Z(n18) );
  CENX1 U1402 ( .A(n1661), .B(a[2]), .Z(n15) );
  CEOX1 U1403 ( .A(a[2]), .B(n1720), .Z(n1457) );
  CENX1 U1404 ( .A(n1712), .B(n1710), .Z(n1200) );
  COND1XL U1405 ( .A(n295), .B(n299), .C(n296), .Z(n294) );
  CND3X1 U1406 ( .A(n1578), .B(n1579), .C(n1580), .Z(n462) );
  CANR1X1 U1407 ( .A(n312), .B(n293), .C(n294), .Z(n292) );
  CANR1X1 U1408 ( .A(n288), .B(n1673), .C(n283), .Z(n281) );
  CNR2X1 U1409 ( .A(n245), .B(n261), .Z(n243) );
  CNR2X1 U1410 ( .A(n791), .B(n800), .Z(n333) );
  CNR2X1 U1411 ( .A(n767), .B(n778), .Z(n322) );
  CNIVX2 U1412 ( .A(n116), .Z(n1746) );
  CIVX2 U1413 ( .A(a[0]), .Z(n6) );
  CANR1XL U1414 ( .A(n365), .B(n1679), .C(n362), .Z(n360) );
  CANR1XL U1415 ( .A(n381), .B(n1681), .C(n378), .Z(n376) );
  CENX1 U1416 ( .A(n297), .B(n179), .Z(product[18]) );
  COND2X1 U1417 ( .A(n36), .B(n1327), .C(n1326), .D(n1658), .Z(n1043) );
  CEOX1 U1418 ( .A(a[24]), .B(n1716), .Z(n1657) );
  COND2X1 U1419 ( .A(n1198), .B(n85), .C(n1197), .D(n82), .Z(n920) );
  COND2X1 U1420 ( .A(n69), .B(n1234), .C(n1233), .D(n66), .Z(n954) );
  CND2X2 U1421 ( .A(n1610), .B(n66), .Z(n69) );
  CIVX2 U1422 ( .A(n1737), .Z(n1735) );
  CIVX2 U1423 ( .A(n1737), .Z(n1734) );
  CIVX2 U1424 ( .A(n39), .Z(n1742) );
  CIVDX1 U1425 ( .A(n89), .Z0(n1562), .Z1(n1563) );
  CIVX2 U1426 ( .A(n30), .Z(n1737) );
  CIVX2 U1427 ( .A(n1711), .Z(n1639) );
  CNIVX1 U1428 ( .A(n909), .Z(n1564) );
  CIVDX1 U1429 ( .A(n3), .Z0(n1565), .Z1(n1566) );
  CIVX1 U1430 ( .A(n1732), .Z(n1727) );
  COND2X1 U1431 ( .A(n77), .B(n1213), .C(n1212), .D(n74), .Z(n934) );
  COND2X1 U1432 ( .A(n97), .B(n1169), .C(n95), .D(n1168), .Z(n893) );
  COND2X1 U1433 ( .A(n97), .B(n1163), .C(n1162), .D(n95), .Z(n887) );
  CAOR1XL U1434 ( .A(n312), .B(n293), .C(n294), .Z(n1571) );
  CNIVX3 U1435 ( .A(n63), .Z(n1711) );
  CENX1 U1436 ( .A(n1713), .B(a[20]), .Z(n89) );
  CAN2X1 U1437 ( .A(n1651), .B(n383), .Z(product[1]) );
  CEOX1 U1438 ( .A(a[26]), .B(n1717), .Z(n1445) );
  CND2X4 U1439 ( .A(n1657), .B(n100), .Z(n102) );
  CFA1XL U1440 ( .A(n997), .B(n1043), .CI(n1019), .CO(n816), .S(n817) );
  COND1X1 U1441 ( .A(n214), .B(n242), .C(n1575), .Z(n1573) );
  COND1X1 U1442 ( .A(n214), .B(n242), .C(n1575), .Z(n213) );
  CEOX1 U1443 ( .A(a[20]), .B(n1714), .Z(n1448) );
  CNR2X2 U1444 ( .A(n513), .B(n538), .Z(n223) );
  CND2XL U1445 ( .A(n1674), .B(n394), .Z(n261) );
  CND2XL U1446 ( .A(n1674), .B(n270), .Z(n175) );
  CND2X2 U1447 ( .A(n89), .B(n1614), .Z(n91) );
  COR2X1 U1448 ( .A(n459), .B(n486), .Z(n1665) );
  COND2X1 U1449 ( .A(n27), .B(n1345), .C(n1653), .D(n1344), .Z(n1060) );
  COND2X1 U1450 ( .A(n44), .B(n1283), .C(n1282), .D(n1654), .Z(n1000) );
  CENX1 U1451 ( .A(n1568), .B(n152), .Z(n1260) );
  CND2X1 U1452 ( .A(n1593), .B(n1594), .Z(n105) );
  CENX4 U1453 ( .A(n1715), .B(a[24]), .Z(n100) );
  CND2XL U1454 ( .A(n263), .B(n1664), .Z(n252) );
  CIVX2 U1455 ( .A(n1569), .Z(n1744) );
  CND2IX2 U1456 ( .B(n1656), .A(n50), .Z(n53) );
  CENX4 U1457 ( .A(n1738), .B(a[10]), .Z(n50) );
  COND2X1 U1458 ( .A(n53), .B(n1275), .C(n1274), .D(n50), .Z(n993) );
  COND2X1 U1459 ( .A(n53), .B(n1259), .C(n1258), .D(n50), .Z(n977) );
  CFA1XL U1460 ( .A(n1041), .B(n1095), .CI(n1067), .CO(n796), .S(n797) );
  COND2X1 U1461 ( .A(n27), .B(n1343), .C(n1653), .D(n1342), .Z(n1058) );
  COND2XL U1462 ( .A(n44), .B(n1281), .C(n1280), .D(n1654), .Z(n998) );
  COND2XL U1463 ( .A(n44), .B(n1282), .C(n1281), .D(n1654), .Z(n999) );
  COND2XL U1464 ( .A(n44), .B(n1294), .C(n1293), .D(n1654), .Z(n1011) );
  COND2XL U1465 ( .A(n44), .B(n1288), .C(n1287), .D(n1654), .Z(n1005) );
  COND2XL U1466 ( .A(n44), .B(n1301), .C(n1300), .D(n1654), .Z(n1018) );
  COND2XL U1467 ( .A(n44), .B(n1742), .C(n1304), .D(n1654), .Z(n861) );
  COND2XL U1468 ( .A(n44), .B(n1285), .C(n1284), .D(n1654), .Z(n1002) );
  COND2XL U1469 ( .A(n44), .B(n1291), .C(n1290), .D(n1654), .Z(n1008) );
  CNR2IXL U1470 ( .B(n1746), .A(n1654), .Z(n1021) );
  COND2XL U1471 ( .A(n44), .B(n1303), .C(n1302), .D(n1654), .Z(n1020) );
  COND2XL U1472 ( .A(n44), .B(n1298), .C(n1297), .D(n1654), .Z(n1015) );
  CEOX2 U1473 ( .A(a[22]), .B(n1715), .Z(n1447) );
  COND2X1 U1474 ( .A(n97), .B(n1168), .C(n95), .D(n1167), .Z(n892) );
  CENXL U1475 ( .A(n1714), .B(n1706), .Z(n1172) );
  CENXL U1476 ( .A(n1661), .B(n1706), .Z(n1412) );
  COND2XL U1477 ( .A(n69), .B(n1223), .C(n1222), .D(n66), .Z(n943) );
  CENXL U1478 ( .A(n1735), .B(n1706), .Z(n1319) );
  CENX2 U1479 ( .A(n1717), .B(a[28]), .Z(n110) );
  CND2X1 U1480 ( .A(n216), .B(n228), .Z(n214) );
  CNR2X1 U1481 ( .A(n234), .B(n239), .Z(n228) );
  CIVXL U1482 ( .A(n312), .Z(n311) );
  CFA1XL U1483 ( .A(n897), .B(n977), .CI(n923), .CO(n452), .S(n453) );
  CFA1XL U1484 ( .A(n985), .B(n1115), .CI(n1031), .CO(n642), .S(n643) );
  COND2X1 U1485 ( .A(n36), .B(n1312), .C(n1311), .D(n1658), .Z(n1028) );
  CNIVX4 U1486 ( .A(n71), .Z(n1712) );
  CHA1X1 U1487 ( .A(n859), .B(n1094), .CO(n788), .S(n789) );
  CFA1X1 U1488 ( .A(n1039), .B(n788), .CI(n1123), .CO(n772), .S(n773) );
  CNR2X1 U1489 ( .A(n322), .B(n327), .Z(n320) );
  CANR1X1 U1490 ( .A(n1665), .B(n213), .C(n210), .Z(n208) );
  CIVDXL U1491 ( .A(n330), .Z0(n329) );
  COND2XL U1492 ( .A(n36), .B(n1324), .C(n1323), .D(n1658), .Z(n1040) );
  COND2XL U1493 ( .A(n36), .B(n1315), .C(n1314), .D(n1658), .Z(n1031) );
  COND2XL U1494 ( .A(n36), .B(n1313), .C(n1312), .D(n1658), .Z(n1029) );
  COND2XL U1495 ( .A(n36), .B(n1325), .C(n1324), .D(n1658), .Z(n1041) );
  CND2X4 U1496 ( .A(n1455), .B(n1658), .Z(n36) );
  CANR1X1 U1497 ( .A(n1663), .B(n1573), .C(n1662), .Z(n199) );
  COND1X1 U1498 ( .A(n280), .B(n292), .C(n281), .Z(n1574) );
  COAN1XL U1499 ( .A(n240), .B(n234), .C(n235), .Z(n1576) );
  CANR1XL U1500 ( .A(n229), .B(n216), .C(n217), .Z(n215) );
  CND2X1 U1501 ( .A(n539), .B(n562), .Z(n235) );
  CNR2X2 U1502 ( .A(n539), .B(n562), .Z(n234) );
  CANR1X2 U1503 ( .A(n257), .B(n1666), .C(n248), .Z(n246) );
  COND1X1 U1504 ( .A(n226), .B(n218), .C(n219), .Z(n217) );
  CND2X1 U1505 ( .A(n1711), .B(a[16]), .Z(n1641) );
  CENXL U1506 ( .A(n1704), .B(n1715), .Z(n1161) );
  COND2XL U1507 ( .A(n97), .B(n1164), .C(n1163), .D(n95), .Z(n888) );
  COND2XL U1508 ( .A(n97), .B(n1165), .C(n1164), .D(n95), .Z(n889) );
  COND2XL U1509 ( .A(n1170), .B(n97), .C(n95), .D(n1169), .Z(n894) );
  CENXL U1510 ( .A(n1745), .B(n1715), .Z(n1170) );
  CENXL U1511 ( .A(n1701), .B(n1715), .Z(n1164) );
  CND2IXL U1512 ( .B(n1746), .A(n1715), .Z(n1171) );
  CENXL U1513 ( .A(n1698), .B(n1715), .Z(n1167) );
  CENXL U1514 ( .A(n1699), .B(n1715), .Z(n1166) );
  CENXL U1515 ( .A(n1702), .B(n1715), .Z(n1163) );
  CENXL U1516 ( .A(n1700), .B(n1715), .Z(n1165) );
  CENXL U1517 ( .A(n1697), .B(n1715), .Z(n1168) );
  CENXL U1518 ( .A(n1703), .B(n1715), .Z(n1162) );
  COND2X1 U1519 ( .A(n18), .B(n1364), .C(n1632), .D(n1363), .Z(n1078) );
  CIVX2 U1520 ( .A(n1583), .Z(n241) );
  CIVX1 U1521 ( .A(n259), .Z(n257) );
  CND2XL U1522 ( .A(n389), .B(n235), .Z(n171) );
  CFA1XL U1523 ( .A(n940), .B(n1050), .CI(n1000), .CO(n476), .S(n477) );
  CENXL U1524 ( .A(n1570), .B(n1706), .Z(n1244) );
  CENXL U1525 ( .A(n1570), .B(n1698), .Z(n1252) );
  CENXL U1526 ( .A(n1570), .B(n1699), .Z(n1251) );
  CENX4 U1527 ( .A(n1570), .B(a[14]), .Z(n66) );
  CNR2X1 U1528 ( .A(n295), .B(n298), .Z(n293) );
  CNR2X2 U1529 ( .A(n707), .B(n722), .Z(n295) );
  CEOX1 U1530 ( .A(n494), .B(n469), .Z(n1577) );
  CEOX1 U1531 ( .A(n1577), .B(n492), .Z(n463) );
  CND2X1 U1532 ( .A(n492), .B(n469), .Z(n1578) );
  CND2X1 U1533 ( .A(n492), .B(n494), .Z(n1579) );
  CND2X1 U1534 ( .A(n469), .B(n494), .Z(n1580) );
  COR2X1 U1535 ( .A(n77), .B(n1205), .Z(n1581) );
  COR2XL U1536 ( .A(n1204), .B(n74), .Z(n1582) );
  CANR1X2 U1537 ( .A(n279), .B(n243), .C(n244), .Z(n1583) );
  CANR1X1 U1538 ( .A(n1574), .B(n243), .C(n244), .Z(n242) );
  COND1X2 U1539 ( .A(n245), .B(n262), .C(n246), .Z(n244) );
  CENXL U1540 ( .A(n1730), .B(n150), .Z(n1343) );
  CIVXL U1541 ( .A(n207), .Z(n205) );
  CNIVX4 U1542 ( .A(n87), .Z(n1714) );
  CND2XL U1543 ( .A(n1665), .B(n212), .Z(n168) );
  CIVX1 U1544 ( .A(n212), .Z(n210) );
  COND1X1 U1545 ( .A(n240), .B(n234), .C(n235), .Z(n229) );
  CND2XL U1546 ( .A(a[28]), .B(n109), .Z(n1585) );
  CND2X1 U1547 ( .A(n1584), .B(n1469), .Z(n1586) );
  CND2X1 U1548 ( .A(n1585), .B(n1586), .Z(n1659) );
  CIVX2 U1549 ( .A(a[28]), .Z(n1584) );
  COR2XL U1550 ( .A(n1263), .B(n50), .Z(n1588) );
  COR2X1 U1551 ( .A(n112), .B(n1142), .Z(n1589) );
  COR2X1 U1552 ( .A(n110), .B(n1141), .Z(n1590) );
  CND2X1 U1553 ( .A(n1589), .B(n1590), .Z(n869) );
  CND2IX2 U1554 ( .B(n1659), .A(n110), .Z(n112) );
  CND2XL U1555 ( .A(n1716), .B(a[26]), .Z(n1593) );
  CND2X1 U1556 ( .A(n1591), .B(n1592), .Z(n1594) );
  CIVXL U1557 ( .A(n1716), .Z(n1591) );
  CIVX2 U1558 ( .A(a[26]), .Z(n1592) );
  COND2XL U1559 ( .A(n107), .B(n1146), .C(n105), .D(n1145), .Z(n872) );
  COND2XL U1560 ( .A(n107), .B(n1148), .C(n105), .D(n1147), .Z(n874) );
  CND2X1 U1561 ( .A(n390), .B(n241), .Z(n1595) );
  CIVX2 U1562 ( .A(n238), .Z(n1596) );
  CND2X1 U1563 ( .A(n1595), .B(n1596), .Z(n1648) );
  CIVXL U1564 ( .A(n239), .Z(n390) );
  CIVXL U1565 ( .A(n240), .Z(n238) );
  CENXL U1566 ( .A(n171), .B(n1648), .Z(product[26]) );
  CIVXL U1567 ( .A(a[14]), .Z(n1597) );
  CIVX2 U1568 ( .A(n1451), .Z(n1609) );
  CENXL U1569 ( .A(n1712), .B(n1709), .Z(n1201) );
  CND2IXL U1570 ( .B(n1746), .A(n1712), .Z(n1216) );
  CENXL U1571 ( .A(n1712), .B(n1705), .Z(n1205) );
  CENXL U1572 ( .A(n1712), .B(n1706), .Z(n1204) );
  CND2X1 U1573 ( .A(n1712), .B(a[18]), .Z(n1646) );
  CIVXL U1574 ( .A(n1083), .Z(n1600) );
  CIVX1 U1575 ( .A(n1600), .Z(n1601) );
  CHA1XL U1576 ( .A(n990), .B(n857), .CO(n736), .S(n737) );
  COND2XL U1577 ( .A(n53), .B(n1258), .C(n1257), .D(n50), .Z(n976) );
  COND2XL U1578 ( .A(n53), .B(n1274), .C(n1273), .D(n50), .Z(n992) );
  COND2XL U1579 ( .A(n53), .B(n1271), .C(n1270), .D(n50), .Z(n989) );
  CNR2IXL U1580 ( .B(n1746), .A(n50), .Z(n997) );
  COND2XL U1581 ( .A(n53), .B(n1278), .C(n1277), .D(n50), .Z(n996) );
  COND2XL U1582 ( .A(n53), .B(n1260), .C(n1259), .D(n50), .Z(n978) );
  COND2XL U1583 ( .A(n53), .B(n1266), .C(n1265), .D(n50), .Z(n984) );
  COND2XL U1584 ( .A(n53), .B(n1261), .C(n1260), .D(n50), .Z(n979) );
  COND2XL U1585 ( .A(n53), .B(n1265), .C(n1264), .D(n50), .Z(n983) );
  COND2XL U1586 ( .A(n53), .B(n1267), .C(n1266), .D(n50), .Z(n985) );
  COND2XL U1587 ( .A(n53), .B(n1567), .C(n1279), .D(n50), .Z(n860) );
  COND2XL U1588 ( .A(n53), .B(n1269), .C(n1268), .D(n50), .Z(n987) );
  COND2XL U1589 ( .A(n53), .B(n1277), .C(n1276), .D(n50), .Z(n995) );
  COND2XL U1590 ( .A(n53), .B(n1276), .C(n1275), .D(n50), .Z(n994) );
  COND2XL U1591 ( .A(n53), .B(n1272), .C(n1271), .D(n50), .Z(n990) );
  CIVX2 U1592 ( .A(n1609), .Z(n1610) );
  CENXL U1593 ( .A(n1745), .B(n1568), .Z(n1278) );
  CND2IXL U1594 ( .B(n1746), .A(n1568), .Z(n1279) );
  CENXL U1595 ( .A(n1568), .B(n1707), .Z(n1266) );
  CENXL U1596 ( .A(n1568), .B(n1705), .Z(n1268) );
  CENXL U1597 ( .A(n1568), .B(n1709), .Z(n1264) );
  CENXL U1598 ( .A(n1568), .B(n151), .Z(n1261) );
  CENXL U1599 ( .A(n1568), .B(n1706), .Z(n1267) );
  CENXL U1600 ( .A(n1568), .B(n1710), .Z(n1263) );
  CENXL U1601 ( .A(n1568), .B(n150), .Z(n1262) );
  CENXL U1602 ( .A(n1568), .B(n1704), .Z(n1269) );
  CIVXL U1603 ( .A(n944), .Z(n1602) );
  CIVX1 U1604 ( .A(n1602), .Z(n1603) );
  CIVX1 U1605 ( .A(n1562), .Z(n1604) );
  CIVXL U1606 ( .A(n261), .Z(n263) );
  CANR1X2 U1607 ( .A(n275), .B(n1674), .C(n268), .Z(n262) );
  CIVX1 U1608 ( .A(n1646), .Z(n1605) );
  CIVX2 U1609 ( .A(n1605), .Z(n1606) );
  CIVX1 U1610 ( .A(n1641), .Z(n1607) );
  CIVX2 U1611 ( .A(n1607), .Z(n1608) );
  CIVXL U1612 ( .A(n1574), .Z(n278) );
  CENXL U1613 ( .A(n1660), .B(n168), .Z(product[29]) );
  CIVX1 U1614 ( .A(n1448), .Z(n1613) );
  CIVX2 U1615 ( .A(n1725), .Z(n1720) );
  CIVX2 U1616 ( .A(n1725), .Z(n1723) );
  CIVX2 U1617 ( .A(n1611), .Z(n1612) );
  CIVX1 U1618 ( .A(n1613), .Z(n1614) );
  CENXL U1619 ( .A(n1683), .B(n220), .Z(product[28]) );
  CENXL U1620 ( .A(n1684), .B(n227), .Z(product[27]) );
  CIVXL U1621 ( .A(n946), .Z(n1615) );
  CIVX2 U1622 ( .A(n1615), .Z(n1616) );
  CENX2 U1623 ( .A(n1743), .B(a[12]), .Z(n58) );
  CIVXL U1624 ( .A(n947), .Z(n1618) );
  CIVX2 U1625 ( .A(n1618), .Z(n1619) );
  CIVXL U1626 ( .A(n945), .Z(n1620) );
  CIVX2 U1627 ( .A(n1620), .Z(n1621) );
  CENXL U1628 ( .A(n1696), .B(n1715), .Z(n1169) );
  CND2X4 U1629 ( .A(n1449), .B(n82), .Z(n85) );
  CEOX1 U1630 ( .A(a[18]), .B(n1713), .Z(n1449) );
  CIVXL U1631 ( .A(n943), .Z(n1622) );
  CIVX2 U1632 ( .A(n1622), .Z(n1623) );
  CIVXL U1633 ( .A(n952), .Z(n1624) );
  CIVX2 U1634 ( .A(n1624), .Z(n1625) );
  CND2X4 U1635 ( .A(n1450), .B(n74), .Z(n77) );
  CEOX1 U1636 ( .A(a[16]), .B(n1712), .Z(n1450) );
  CIVX2 U1637 ( .A(a[8]), .Z(n1629) );
  CIVX4 U1638 ( .A(n1629), .Z(n1630) );
  CENX1 U1639 ( .A(n1661), .B(a[2]), .Z(n1631) );
  CENX1 U1640 ( .A(n1661), .B(a[2]), .Z(n1632) );
  CNR2XL U1641 ( .A(n18), .B(n1381), .Z(n1633) );
  CNR2XL U1642 ( .A(n1631), .B(n1380), .Z(n1634) );
  COR2X1 U1643 ( .A(n1633), .B(n1634), .Z(n1095) );
  CIVX1 U1644 ( .A(n1723), .Z(n1635) );
  CIVX2 U1645 ( .A(a[4]), .Z(n1636) );
  COND2XL U1646 ( .A(n27), .B(n1347), .C(n1653), .D(n1346), .Z(n1062) );
  COND2XL U1647 ( .A(n27), .B(n1338), .C(n1653), .D(n1337), .Z(n1053) );
  COND2XL U1648 ( .A(n27), .B(n1355), .C(n1653), .D(n1354), .Z(n1070) );
  COND2XL U1649 ( .A(n27), .B(n1350), .C(n1653), .D(n1349), .Z(n1065) );
  COND2XL U1650 ( .A(n27), .B(n1340), .C(n1653), .D(n1339), .Z(n1055) );
  COND2XL U1651 ( .A(n27), .B(n1335), .C(n1653), .D(n1334), .Z(n1050) );
  COND2XL U1652 ( .A(n27), .B(n1354), .C(n1653), .D(n1353), .Z(n1069) );
  COND2XL U1653 ( .A(n27), .B(n1356), .C(n1653), .D(n1355), .Z(n1071) );
  COND2XL U1654 ( .A(n27), .B(n1334), .C(n1653), .D(n1333), .Z(n1049) );
  COND2XL U1655 ( .A(n27), .B(n1333), .C(n1653), .D(n1332), .Z(n1048) );
  CNR2IX1 U1656 ( .B(n1746), .A(n1653), .Z(n1075) );
  COND2XL U1657 ( .A(n27), .B(n1351), .C(n1653), .D(n1350), .Z(n1066) );
  COND2XL U1658 ( .A(n27), .B(n1342), .C(n1653), .D(n1341), .Z(n1057) );
  COND2XL U1659 ( .A(n27), .B(n1339), .C(n1653), .D(n1338), .Z(n1054) );
  COND2XL U1660 ( .A(n27), .B(n1341), .C(n1653), .D(n1340), .Z(n1056) );
  COND2XL U1661 ( .A(n27), .B(n1353), .C(n1653), .D(n1352), .Z(n1068) );
  COND2XL U1662 ( .A(n27), .B(n1732), .C(n1360), .D(n1653), .Z(n863) );
  COND2XL U1663 ( .A(n27), .B(n1336), .C(n1653), .D(n1335), .Z(n1051) );
  COND2XL U1664 ( .A(n27), .B(n1357), .C(n1653), .D(n1356), .Z(n1072) );
  COND2XL U1665 ( .A(n27), .B(n1359), .C(n1653), .D(n1358), .Z(n1074) );
  COND2XL U1666 ( .A(n27), .B(n1358), .C(n1653), .D(n1357), .Z(n1073) );
  CENXL U1667 ( .A(n1711), .B(n150), .Z(n1218) );
  CND2IXL U1668 ( .B(n1746), .A(n1711), .Z(n1235) );
  CENXL U1669 ( .A(n1711), .B(n1696), .Z(n1233) );
  CND2X2 U1670 ( .A(n1639), .B(n1640), .Z(n1642) );
  CND2X4 U1671 ( .A(n1608), .B(n1642), .Z(n74) );
  CIVX2 U1672 ( .A(a[16]), .Z(n1640) );
  COND2XL U1673 ( .A(n77), .B(n1201), .C(n1200), .D(n74), .Z(n922) );
  COND2XL U1674 ( .A(n77), .B(n1644), .C(n74), .D(n1216), .Z(n857) );
  COND2XL U1675 ( .A(n1215), .B(n77), .C(n1214), .D(n74), .Z(n936) );
  CIVXL U1676 ( .A(n234), .Z(n389) );
  COND2X1 U1677 ( .A(n85), .B(n1194), .C(n1193), .D(n82), .Z(n916) );
  CIVXL U1678 ( .A(a[18]), .Z(n1645) );
  CNR2IX1 U1679 ( .B(n1746), .A(n82), .Z(n921) );
  CIVXL U1680 ( .A(n1713), .Z(n1474) );
  CIVXL U1681 ( .A(n1715), .Z(n1472) );
  CIVXL U1682 ( .A(n264), .Z(n1643) );
  CIVXL U1683 ( .A(n262), .Z(n264) );
  CND2X4 U1684 ( .A(n1606), .B(n1647), .Z(n82) );
  CIVXL U1685 ( .A(n1712), .Z(n1644) );
  COND2XL U1686 ( .A(n85), .B(n1186), .C(n1185), .D(n82), .Z(n908) );
  COND2XL U1687 ( .A(n85), .B(n1189), .C(n1188), .D(n82), .Z(n911) );
  CEOX2 U1688 ( .A(a[12]), .B(n1626), .Z(n1452) );
  CIVX2 U1689 ( .A(n1742), .Z(n1738) );
  CENX1 U1690 ( .A(n1627), .B(n1708), .Z(n1242) );
  CENX1 U1691 ( .A(n1628), .B(n1710), .Z(n1240) );
  CENX1 U1692 ( .A(n1628), .B(n1709), .Z(n1241) );
  CENX1 U1693 ( .A(n1746), .B(n1627), .Z(n1255) );
  CNIVX2 U1694 ( .A(n136), .Z(n1704) );
  CANR1X1 U1695 ( .A(n1670), .B(n321), .C(n316), .Z(n314) );
  CND2IXL U1696 ( .B(n1746), .A(n1627), .Z(n1256) );
  COND2XL U1697 ( .A(n69), .B(n1220), .C(n1219), .D(n66), .Z(n940) );
  CNIVX2 U1698 ( .A(n116), .Z(n1745) );
  CIVX2 U1699 ( .A(n12), .Z(n1725) );
  CND2XL U1700 ( .A(n397), .B(n296), .Z(n179) );
  CNR2X1 U1701 ( .A(n739), .B(n752), .Z(n305) );
  CND2XL U1702 ( .A(n430), .B(n415), .Z(n198) );
  CENX1 U1703 ( .A(n191), .B(n365), .Z(product[6]) );
  CND2XL U1704 ( .A(n412), .B(n375), .Z(n194) );
  COND2XL U1705 ( .A(n44), .B(n1287), .C(n1286), .D(n1654), .Z(n1004) );
  CNIVX4 U1706 ( .A(n1728), .Z(n1682) );
  CND2X4 U1707 ( .A(n1458), .B(n6), .Z(n9) );
  CENX1 U1708 ( .A(a[4]), .B(n1731), .Z(n1652) );
  CNIVX1 U1709 ( .A(n140), .Z(n1706) );
  CNIVX2 U1710 ( .A(n132), .Z(n1702) );
  CNIVX1 U1711 ( .A(n144), .Z(n1708) );
  CNIVX1 U1712 ( .A(n146), .Z(n1709) );
  CENXL U1713 ( .A(n1686), .B(n208), .Z(product[30]) );
  CND2XL U1714 ( .A(n390), .B(n240), .Z(n172) );
  CNR2IXL U1715 ( .B(n228), .A(n223), .Z(n221) );
  CAN2XL U1716 ( .A(n1667), .B(n1665), .Z(n1663) );
  CIVX1 U1717 ( .A(n270), .Z(n268) );
  CANR1X1 U1718 ( .A(n308), .B(n1671), .C(n301), .Z(n299) );
  CIVX1 U1719 ( .A(n303), .Z(n301) );
  CND2XL U1720 ( .A(n1670), .B(n318), .Z(n182) );
  CEOXL U1721 ( .A(n182), .B(n319), .Z(product[15]) );
  CEOXL U1722 ( .A(n177), .B(n286), .Z(product[20]) );
  CND2XL U1723 ( .A(n1673), .B(n285), .Z(n177) );
  CEOXL U1724 ( .A(n176), .B(n278), .Z(product[21]) );
  CND2XL U1725 ( .A(n394), .B(n273), .Z(n176) );
  CEOXL U1726 ( .A(n181), .B(n311), .Z(product[16]) );
  CND2XL U1727 ( .A(n399), .B(n306), .Z(n181) );
  CEOXL U1728 ( .A(n183), .B(n324), .Z(product[14]) );
  CND2XL U1729 ( .A(n1672), .B(n290), .Z(n178) );
  CND2XL U1730 ( .A(n1671), .B(n399), .Z(n298) );
  CND2XL U1731 ( .A(n404), .B(n337), .Z(n186) );
  CEOXL U1732 ( .A(n186), .B(n338), .Z(product[11]) );
  CEOXL U1733 ( .A(n346), .B(n187), .Z(product[10]) );
  CND2XL U1734 ( .A(n1676), .B(n345), .Z(n187) );
  CND2XL U1735 ( .A(n402), .B(n328), .Z(n184) );
  CND2XL U1736 ( .A(n1677), .B(n356), .Z(n189) );
  CND2XL U1737 ( .A(n1675), .B(n350), .Z(n188) );
  CND2XL U1738 ( .A(n767), .B(n778), .Z(n323) );
  CND2XL U1739 ( .A(n707), .B(n722), .Z(n296) );
  CENX1 U1740 ( .A(n1649), .B(n653), .Z(n651) );
  CENX1 U1741 ( .A(n655), .B(n672), .Z(n1649) );
  CENXL U1742 ( .A(n1685), .B(n199), .Z(product[31]) );
  CANR1X1 U1743 ( .A(n373), .B(n1680), .C(n370), .Z(n368) );
  CND2IXL U1744 ( .B(n366), .A(n367), .Z(n192) );
  CND2IXL U1745 ( .B(n358), .A(n359), .Z(n190) );
  CND2XL U1746 ( .A(n1679), .B(n364), .Z(n191) );
  CND2XL U1747 ( .A(n791), .B(n800), .Z(n334) );
  CND2XL U1748 ( .A(n1681), .B(n380), .Z(n195) );
  CEOXL U1749 ( .A(n376), .B(n194), .Z(product[3]) );
  CND2XL U1750 ( .A(n849), .B(n864), .Z(n375) );
  CEN3X1 U1751 ( .A(n434), .B(n1650), .C(n432), .Z(n415) );
  CEN3X2 U1752 ( .A(n436), .B(n418), .C(n417), .Z(n1650) );
  CEO3X1 U1753 ( .A(n452), .B(n450), .C(n448), .Z(n422) );
  COR2XL U1754 ( .A(n1136), .B(n865), .Z(n1651) );
  COND2XL U1755 ( .A(n18), .B(n1387), .C(n1632), .D(n1386), .Z(n1101) );
  CNR2IXL U1756 ( .B(n1746), .A(n1631), .Z(n1105) );
  CNR2IXL U1757 ( .B(n1746), .A(n100), .Z(n885) );
  COND2XL U1758 ( .A(n97), .B(n1162), .C(n1161), .D(n95), .Z(n886) );
  CNIVX4 U1759 ( .A(n3), .Z(n1661) );
  CEOX2 U1760 ( .A(a[0]), .B(n1718), .Z(n1458) );
  CND2X4 U1761 ( .A(n1452), .B(n58), .Z(n61) );
  CENX2 U1762 ( .A(n1714), .B(a[22]), .Z(n95) );
  CENX4 U1763 ( .A(n1734), .B(n1630), .Z(n1654) );
  CND2IX4 U1764 ( .B(n1655), .A(n1654), .Z(n44) );
  CENX1 U1765 ( .A(n1630), .B(n1741), .Z(n1655) );
  CENX4 U1766 ( .A(n1682), .B(a[6]), .Z(n1658) );
  CNIVX2 U1767 ( .A(n142), .Z(n1707) );
  CND2XL U1768 ( .A(n1443), .B(n114), .Z(n115) );
  CIVXL U1769 ( .A(n109), .Z(n1469) );
  COND1XL U1770 ( .A(n214), .B(n1583), .C(n215), .Z(n1660) );
  COND1X1 U1771 ( .A(n330), .B(n313), .C(n314), .Z(n312) );
  CENX1 U1772 ( .A(n241), .B(n172), .Z(product[25]) );
  CANR1XL U1773 ( .A(n228), .B(n241), .C(n229), .Z(n227) );
  CANR1XL U1774 ( .A(n221), .B(n241), .C(n222), .Z(n220) );
  CANR1XL U1775 ( .A(n1664), .B(n264), .C(n257), .Z(n253) );
  CNR2X1 U1776 ( .A(n218), .B(n223), .Z(n216) );
  CENX1 U1777 ( .A(n260), .B(n174), .Z(product[23]) );
  COND1XL U1778 ( .A(n261), .B(n278), .C(n1643), .Z(n260) );
  CENX1 U1779 ( .A(n251), .B(n173), .Z(product[24]) );
  COND1XL U1780 ( .A(n252), .B(n278), .C(n253), .Z(n251) );
  COND1XL U1781 ( .A(n223), .B(n1576), .C(n226), .Z(n222) );
  CAOR1X1 U1782 ( .A(n210), .B(n1667), .C(n205), .Z(n1662) );
  CND2X1 U1783 ( .A(n320), .B(n1670), .Z(n313) );
  CNR2X1 U1784 ( .A(n487), .B(n512), .Z(n218) );
  COND1X1 U1785 ( .A(n280), .B(n292), .C(n281), .Z(n279) );
  CND2X1 U1786 ( .A(n1673), .B(n1672), .Z(n280) );
  CENX1 U1787 ( .A(n271), .B(n175), .Z(product[22]) );
  COND1XL U1788 ( .A(n272), .B(n278), .C(n273), .Z(n271) );
  CENX1 U1789 ( .A(n304), .B(n180), .Z(product[17]) );
  CND2X1 U1790 ( .A(n1671), .B(n303), .Z(n180) );
  COND1XL U1791 ( .A(n305), .B(n311), .C(n306), .Z(n304) );
  CENX1 U1792 ( .A(n1571), .B(n178), .Z(product[19]) );
  CANR1XL U1793 ( .A(n1672), .B(n1571), .C(n288), .Z(n286) );
  CND2X1 U1794 ( .A(n401), .B(n323), .Z(n183) );
  CANR1XL U1795 ( .A(n402), .B(n329), .C(n326), .Z(n324) );
  COR2X1 U1796 ( .A(n609), .B(n630), .Z(n1664) );
  CND2X1 U1797 ( .A(n563), .B(n586), .Z(n240) );
  COR2X1 U1798 ( .A(n587), .B(n608), .Z(n1666) );
  CND2X1 U1799 ( .A(n459), .B(n486), .Z(n212) );
  CND2X1 U1800 ( .A(n513), .B(n538), .Z(n226) );
  COR2X1 U1801 ( .A(n431), .B(n458), .Z(n1667) );
  CND2X1 U1802 ( .A(n487), .B(n512), .Z(n219) );
  CND2X1 U1803 ( .A(n609), .B(n630), .Z(n259) );
  CND2X1 U1804 ( .A(n587), .B(n608), .Z(n250) );
  CND2X1 U1805 ( .A(n431), .B(n458), .Z(n207) );
  CENX1 U1806 ( .A(n1668), .B(n489), .Z(n487) );
  CENX1 U1807 ( .A(n514), .B(n491), .Z(n1668) );
  CENX1 U1808 ( .A(n1669), .B(n589), .Z(n587) );
  CENX1 U1809 ( .A(n610), .B(n591), .Z(n1669) );
  COND1XL U1810 ( .A(n352), .B(n340), .C(n341), .Z(n339) );
  CND2X1 U1811 ( .A(n1676), .B(n1675), .Z(n340) );
  CANR1XL U1812 ( .A(n348), .B(n1676), .C(n343), .Z(n341) );
  CANR1X1 U1813 ( .A(n331), .B(n339), .C(n332), .Z(n330) );
  CNR2X1 U1814 ( .A(n333), .B(n336), .Z(n331) );
  COND1XL U1815 ( .A(n337), .B(n333), .C(n334), .Z(n332) );
  CENX1 U1816 ( .A(n189), .B(n357), .Z(product[8]) );
  CENX1 U1817 ( .A(n188), .B(n351), .Z(product[9]) );
  CENX1 U1818 ( .A(n335), .B(n185), .Z(product[12]) );
  CND2X1 U1819 ( .A(n403), .B(n334), .Z(n185) );
  COND1XL U1820 ( .A(n336), .B(n338), .C(n337), .Z(n335) );
  CENX1 U1821 ( .A(n329), .B(n184), .Z(product[13]) );
  CNR2X1 U1822 ( .A(n651), .B(n670), .Z(n272) );
  COR2X1 U1823 ( .A(n753), .B(n766), .Z(n1670) );
  CANR1XL U1824 ( .A(n1675), .B(n351), .C(n348), .Z(n346) );
  COR2X1 U1825 ( .A(n723), .B(n738), .Z(n1671) );
  COR2X1 U1826 ( .A(n689), .B(n706), .Z(n1672) );
  CND2X1 U1827 ( .A(n651), .B(n670), .Z(n273) );
  CND2X1 U1828 ( .A(n739), .B(n752), .Z(n306) );
  COR2X1 U1829 ( .A(n671), .B(n688), .Z(n1673) );
  COR2X1 U1830 ( .A(n631), .B(n650), .Z(n1674) );
  CND2X1 U1831 ( .A(n689), .B(n706), .Z(n290) );
  CND2X1 U1832 ( .A(n631), .B(n650), .Z(n270) );
  CND2X1 U1833 ( .A(n723), .B(n738), .Z(n303) );
  CND2X1 U1834 ( .A(n671), .B(n688), .Z(n285) );
  CND2X1 U1835 ( .A(n753), .B(n766), .Z(n318) );
  COND1XL U1836 ( .A(n376), .B(n374), .C(n375), .Z(n373) );
  COND1XL U1837 ( .A(n368), .B(n366), .C(n367), .Z(n365) );
  CND3XL U1838 ( .A(n1687), .B(n1688), .C(n1689), .Z(n650) );
  CNR2X1 U1839 ( .A(n801), .B(n810), .Z(n336) );
  CNR2X1 U1840 ( .A(n779), .B(n790), .Z(n327) );
  CND2X1 U1841 ( .A(n779), .B(n790), .Z(n328) );
  COR2X1 U1842 ( .A(n819), .B(n826), .Z(n1675) );
  COR2X1 U1843 ( .A(n811), .B(n818), .Z(n1676) );
  CND2X1 U1844 ( .A(n801), .B(n810), .Z(n337) );
  CND2X1 U1845 ( .A(n819), .B(n826), .Z(n350) );
  CND2X1 U1846 ( .A(n811), .B(n818), .Z(n345) );
  CND2X1 U1847 ( .A(n827), .B(n832), .Z(n356) );
  COR2X1 U1848 ( .A(n827), .B(n832), .Z(n1677) );
  COR2X1 U1849 ( .A(n430), .B(n415), .Z(n1678) );
  CENX1 U1850 ( .A(n195), .B(n381), .Z(product[2]) );
  CENX1 U1851 ( .A(n193), .B(n373), .Z(product[4]) );
  CND2X1 U1852 ( .A(n1680), .B(n372), .Z(n193) );
  CNR2X1 U1853 ( .A(n833), .B(n838), .Z(n358) );
  CNR2X1 U1854 ( .A(n849), .B(n864), .Z(n374) );
  CNR2X1 U1855 ( .A(n843), .B(n846), .Z(n366) );
  CND2X1 U1856 ( .A(n833), .B(n838), .Z(n359) );
  CND2X1 U1857 ( .A(n1136), .B(n865), .Z(n383) );
  CND2X1 U1858 ( .A(n847), .B(n848), .Z(n372) );
  CND2X1 U1859 ( .A(n839), .B(n842), .Z(n364) );
  CND2X1 U1860 ( .A(n1135), .B(n1105), .Z(n380) );
  COR2X1 U1861 ( .A(n839), .B(n842), .Z(n1679) );
  CND2X1 U1862 ( .A(n843), .B(n846), .Z(n367) );
  COR2X1 U1863 ( .A(n847), .B(n848), .Z(n1680) );
  COR2X1 U1864 ( .A(n1135), .B(n1105), .Z(n1681) );
  CENX1 U1865 ( .A(n1739), .B(n1707), .Z(n1291) );
  CENX1 U1866 ( .A(n1570), .B(n1701), .Z(n1249) );
  CENX1 U1867 ( .A(n1739), .B(n1706), .Z(n1292) );
  CENX1 U1868 ( .A(n1570), .B(n1704), .Z(n1246) );
  CENX1 U1869 ( .A(n1700), .B(n1717), .Z(n1145) );
  CENX1 U1870 ( .A(n1745), .B(n1718), .Z(n1423) );
  CENX1 U1871 ( .A(n1729), .B(n1707), .Z(n1347) );
  CENX1 U1872 ( .A(n1730), .B(n1710), .Z(n1344) );
  CENX1 U1873 ( .A(n1729), .B(n1706), .Z(n1348) );
  CENX1 U1874 ( .A(n1661), .B(n1698), .Z(n1420) );
  CENX1 U1875 ( .A(n1661), .B(n1700), .Z(n1418) );
  CENX1 U1876 ( .A(n1661), .B(n1701), .Z(n1417) );
  CENX1 U1877 ( .A(n1682), .B(n1704), .Z(n1350) );
  CENX1 U1878 ( .A(n1661), .B(n1704), .Z(n1414) );
  CNR2IX1 U1879 ( .B(n1746), .A(n105), .Z(n877) );
  CIVX2 U1880 ( .A(n1565), .Z(n1718) );
  CENX1 U1881 ( .A(n1713), .B(n1708), .Z(n1185) );
  CIVX2 U1882 ( .A(n1567), .Z(n1743) );
  CENX1 U1883 ( .A(n1702), .B(n1716), .Z(n1152) );
  CENX1 U1884 ( .A(n1722), .B(n1698), .Z(n1387) );
  CENX1 U1885 ( .A(n1722), .B(n1699), .Z(n1386) );
  CENX1 U1886 ( .A(n1739), .B(n1701), .Z(n1297) );
  CENX1 U1887 ( .A(n1739), .B(n1700), .Z(n1298) );
  CENX1 U1888 ( .A(n1740), .B(n1699), .Z(n1299) );
  CENX1 U1889 ( .A(n1740), .B(n1702), .Z(n1296) );
  CENX1 U1890 ( .A(n1735), .B(n1708), .Z(n1317) );
  CENX1 U1891 ( .A(n1735), .B(n1710), .Z(n1315) );
  CENX1 U1892 ( .A(n1735), .B(n1709), .Z(n1316) );
  CENX1 U1893 ( .A(n1713), .B(n1697), .Z(n1196) );
  CENX1 U1894 ( .A(n1714), .B(n1702), .Z(n1176) );
  CENX1 U1895 ( .A(n1713), .B(n1700), .Z(n1193) );
  CENX1 U1896 ( .A(n1740), .B(n1709), .Z(n1289) );
  CENX1 U1897 ( .A(n1741), .B(n1704), .Z(n1294) );
  CENX1 U1898 ( .A(n1735), .B(n1701), .Z(n1324) );
  CENX1 U1899 ( .A(n1740), .B(n1703), .Z(n1295) );
  CENX1 U1900 ( .A(n1714), .B(n1699), .Z(n1179) );
  CENX1 U1901 ( .A(n1714), .B(n1700), .Z(n1178) );
  CENX1 U1902 ( .A(n1713), .B(n1702), .Z(n1191) );
  CENX1 U1903 ( .A(n1713), .B(n1701), .Z(n1192) );
  CENX1 U1904 ( .A(n1735), .B(n1704), .Z(n1321) );
  CENX1 U1905 ( .A(n1696), .B(n1714), .Z(n1182) );
  CENX1 U1906 ( .A(n1713), .B(n1698), .Z(n1195) );
  CENX1 U1907 ( .A(n1739), .B(n1708), .Z(n1290) );
  CENX1 U1908 ( .A(n1714), .B(n1701), .Z(n1177) );
  CENX1 U1909 ( .A(n1713), .B(n1704), .Z(n1189) );
  CENX1 U1910 ( .A(n1713), .B(n1699), .Z(n1194) );
  CENX1 U1911 ( .A(n1714), .B(n1703), .Z(n1175) );
  CENX1 U1912 ( .A(n1740), .B(n1710), .Z(n1288) );
  CENX1 U1913 ( .A(n1697), .B(n1714), .Z(n1181) );
  CENX1 U1914 ( .A(n1698), .B(n1714), .Z(n1180) );
  CENX1 U1915 ( .A(n1714), .B(n1705), .Z(n1173) );
  CENX1 U1916 ( .A(n1714), .B(n1704), .Z(n1174) );
  CENX1 U1917 ( .A(n1713), .B(n1707), .Z(n1186) );
  CENX1 U1918 ( .A(n1713), .B(n1706), .Z(n1187) );
  CENX1 U1919 ( .A(n1566), .B(n1702), .Z(n1416) );
  CENX1 U1920 ( .A(n1724), .B(n1709), .Z(n1376) );
  CENX1 U1921 ( .A(n1727), .B(n1698), .Z(n1356) );
  CENX1 U1922 ( .A(n1729), .B(n1708), .Z(n1346) );
  CENX1 U1923 ( .A(n1727), .B(n1697), .Z(n1357) );
  CENX1 U1924 ( .A(n1729), .B(n1709), .Z(n1345) );
  CENX1 U1925 ( .A(n1661), .B(n1696), .Z(n1422) );
  CENX1 U1926 ( .A(n1661), .B(n1697), .Z(n1421) );
  CENX1 U1927 ( .A(n1661), .B(n1699), .Z(n1419) );
  CENX1 U1928 ( .A(n1727), .B(n1696), .Z(n1358) );
  CENX1 U1929 ( .A(n1718), .B(n1707), .Z(n1411) );
  CENX1 U1930 ( .A(n1718), .B(n1708), .Z(n1410) );
  CENX1 U1931 ( .A(n1697), .B(n1716), .Z(n1157) );
  CENX1 U1932 ( .A(n1696), .B(n1716), .Z(n1158) );
  CENX1 U1933 ( .A(n1724), .B(n1708), .Z(n1377) );
  CENX1 U1934 ( .A(n1718), .B(n1710), .Z(n1408) );
  CENX1 U1935 ( .A(n1718), .B(n1709), .Z(n1409) );
  CENX1 U1936 ( .A(n1699), .B(n1716), .Z(n1155) );
  CENX1 U1937 ( .A(n1698), .B(n1716), .Z(n1156) );
  CENX1 U1938 ( .A(n1698), .B(n1717), .Z(n1147) );
  CENX1 U1939 ( .A(n1701), .B(n1716), .Z(n1153) );
  CENX1 U1940 ( .A(n1700), .B(n1716), .Z(n1154) );
  CENX1 U1941 ( .A(n1699), .B(n1717), .Z(n1146) );
  CENX1 U1942 ( .A(n1735), .B(n1702), .Z(n1323) );
  CENX1 U1943 ( .A(n1734), .B(n1700), .Z(n1325) );
  CENX1 U1944 ( .A(n1734), .B(n1698), .Z(n1327) );
  CENX1 U1945 ( .A(n1733), .B(n1707), .Z(n1318) );
  CENX1 U1946 ( .A(n1735), .B(n1703), .Z(n1322) );
  CENX1 U1947 ( .A(n1724), .B(n1707), .Z(n1378) );
  CENX1 U1948 ( .A(n1721), .B(n1706), .Z(n1379) );
  CENX1 U1949 ( .A(n1724), .B(n1710), .Z(n1375) );
  CENX1 U1950 ( .A(n1745), .B(n1741), .Z(n1303) );
  CENX1 U1951 ( .A(n1745), .B(n1713), .Z(n1198) );
  CENX1 U1952 ( .A(n1745), .B(n1714), .Z(n1183) );
  CENX1 U1953 ( .A(n1745), .B(n1716), .Z(n1159) );
  CENX1 U1954 ( .A(n1745), .B(n1717), .Z(n1150) );
  CENX1 U1955 ( .A(n1734), .B(n1697), .Z(n1328) );
  CENX1 U1956 ( .A(n1735), .B(n1696), .Z(n1329) );
  CENX1 U1957 ( .A(n1745), .B(n1731), .Z(n1359) );
  CENX1 U1958 ( .A(n1722), .B(n1697), .Z(n1388) );
  CENX1 U1959 ( .A(n1722), .B(n1700), .Z(n1385) );
  CENX1 U1960 ( .A(n1719), .B(n1696), .Z(n1389) );
  CENX1 U1961 ( .A(n1721), .B(n1701), .Z(n1384) );
  CENX1 U1962 ( .A(n1721), .B(n1702), .Z(n1383) );
  CENX1 U1963 ( .A(n1745), .B(n1719), .Z(n1390) );
  CNR2IX1 U1964 ( .B(n1746), .A(n1617), .Z(n975) );
  CNR2IX1 U1965 ( .B(n1746), .A(n114), .Z(n867) );
  CNR2IX1 U1966 ( .B(n1746), .A(n1563), .Z(n907) );
  CNR2IX1 U1967 ( .B(n1746), .A(n95), .Z(n895) );
  CNR2IX1 U1968 ( .B(n1746), .A(n110), .Z(n871) );
  CEOX1 U1969 ( .A(n872), .B(n886), .Z(n429) );
  CNR2IX1 U1970 ( .B(n1746), .A(n6), .Z(product[0]) );
  CENX1 U1971 ( .A(n1735), .B(b[25]), .Z(n1305) );
  CENX1 U1972 ( .A(n1721), .B(b[29]), .Z(n1361) );
  CENX1 U1973 ( .A(n1661), .B(n152), .Z(n1405) );
  CENX1 U1974 ( .A(n1724), .B(n151), .Z(n1373) );
  CENX1 U1975 ( .A(n1727), .B(n157), .Z(n1336) );
  CENX1 U1976 ( .A(n1727), .B(n156), .Z(n1337) );
  CENX1 U1977 ( .A(n109), .B(a[30]), .Z(n114) );
  CENX1 U1978 ( .A(n1661), .B(b[31]), .Z(n1392) );
  CENX1 U1979 ( .A(n1727), .B(b[27]), .Z(n1332) );
  CENX1 U1980 ( .A(n1733), .B(n157), .Z(n1307) );
  CENX1 U1981 ( .A(n1733), .B(b[24]), .Z(n1306) );
  CENX1 U1982 ( .A(n1739), .B(n154), .Z(n1283) );
  CENX1 U1983 ( .A(n1745), .B(n113), .Z(n1138) );
  CENX1 U1984 ( .A(n1696), .B(n113), .Z(n1137) );
  CENX1 U1985 ( .A(n1698), .B(n109), .Z(n1140) );
  CENX1 U1986 ( .A(n1740), .B(n151), .Z(n1286) );
  CENX1 U1987 ( .A(n1740), .B(n150), .Z(n1287) );
  CENX1 U1988 ( .A(n1739), .B(n152), .Z(n1285) );
  CENX1 U1989 ( .A(n1735), .B(n150), .Z(n1314) );
  CENX1 U1990 ( .A(n1735), .B(n154), .Z(n1310) );
  CENX1 U1991 ( .A(n1627), .B(n150), .Z(n1239) );
  CENX1 U1992 ( .A(n1739), .B(n156), .Z(n1281) );
  CENX1 U1993 ( .A(n1628), .B(n151), .Z(n1238) );
  CENX1 U1994 ( .A(n1628), .B(n152), .Z(n1237) );
  CENX1 U1995 ( .A(n1566), .B(n153), .Z(n1404) );
  CENX1 U1996 ( .A(n1566), .B(n157), .Z(n1400) );
  CENX1 U1997 ( .A(n1727), .B(n154), .Z(n1339) );
  CENX1 U1998 ( .A(n1727), .B(n155), .Z(n1338) );
  CENX1 U1999 ( .A(n1566), .B(b[24]), .Z(n1399) );
  CENX1 U2000 ( .A(n1566), .B(b[25]), .Z(n1398) );
  CENX1 U2001 ( .A(n1720), .B(n157), .Z(n1367) );
  CENX1 U2002 ( .A(n1566), .B(n156), .Z(n1401) );
  CENX1 U2003 ( .A(n1723), .B(n152), .Z(n1372) );
  CENX1 U2004 ( .A(n1566), .B(n154), .Z(n1403) );
  CENX1 U2005 ( .A(n1566), .B(n155), .Z(n1402) );
  CENX1 U2006 ( .A(n1720), .B(b[24]), .Z(n1366) );
  CENX1 U2007 ( .A(n1566), .B(b[27]), .Z(n1396) );
  CENX1 U2008 ( .A(n1566), .B(b[26]), .Z(n1397) );
  CENX1 U2009 ( .A(n1566), .B(b[28]), .Z(n1395) );
  CENX1 U2010 ( .A(n1718), .B(n151), .Z(n1406) );
  CENX1 U2011 ( .A(n1718), .B(n150), .Z(n1407) );
  CENX1 U2012 ( .A(n1730), .B(b[24]), .Z(n1335) );
  CENX1 U2013 ( .A(n1727), .B(b[25]), .Z(n1334) );
  CENX1 U2014 ( .A(n1727), .B(b[26]), .Z(n1333) );
  CENX1 U2015 ( .A(n1566), .B(b[29]), .Z(n1394) );
  CENX1 U2016 ( .A(n1566), .B(b[30]), .Z(n1393) );
  CENX1 U2017 ( .A(n1720), .B(n156), .Z(n1368) );
  CENX1 U2018 ( .A(n1720), .B(b[25]), .Z(n1365) );
  CENX1 U2019 ( .A(n1721), .B(n154), .Z(n1370) );
  CENX1 U2020 ( .A(n1740), .B(n157), .Z(n1280) );
  CENX1 U2021 ( .A(n1745), .B(n109), .Z(n1143) );
  CENX1 U2022 ( .A(n1719), .B(b[26]), .Z(n1364) );
  CENX1 U2023 ( .A(n1721), .B(n155), .Z(n1369) );
  CENX1 U2024 ( .A(n1719), .B(b[27]), .Z(n1363) );
  CENX1 U2025 ( .A(n1719), .B(b[28]), .Z(n1362) );
  CND2X1 U2026 ( .A(n1445), .B(n105), .Z(n107) );
  CNIVX3 U2027 ( .A(n93), .Z(n1715) );
  CND2X2 U2028 ( .A(n95), .B(n1447), .Z(n97) );
  CEOX1 U2029 ( .A(a[30]), .B(n113), .Z(n1443) );
  CIVX1 U2030 ( .A(n1742), .Z(n1739) );
  CND2XL U2031 ( .A(n1666), .B(n250), .Z(n173) );
  CND2XL U2032 ( .A(n1664), .B(n259), .Z(n174) );
  CIVXL U2033 ( .A(n339), .Z(n338) );
  CFA1XL U2034 ( .A(n1021), .B(n1129), .CI(n1045), .CO(n830), .S(n831) );
  CAN2XL U2035 ( .A(n387), .B(n219), .Z(n1683) );
  CAN2XL U2036 ( .A(n388), .B(n226), .Z(n1684) );
  CAN2X1 U2037 ( .A(n1678), .B(n198), .Z(n1685) );
  CAN2XL U2038 ( .A(n1667), .B(n207), .Z(n1686) );
  CFA1X1 U2039 ( .A(n954), .B(n1092), .CI(n1038), .CO(n760), .S(n761) );
  CENX1 U2040 ( .A(n1730), .B(n151), .Z(n1342) );
  CENX1 U2041 ( .A(n1740), .B(n155), .Z(n1282) );
  CENX1 U2042 ( .A(n1726), .B(n1702), .Z(n1352) );
  CENX1 U2043 ( .A(n1726), .B(n1699), .Z(n1355) );
  CENX1 U2044 ( .A(n1726), .B(n1700), .Z(n1354) );
  CENX1 U2045 ( .A(n1726), .B(n1701), .Z(n1353) );
  CIVX1 U2046 ( .A(n1742), .Z(n1741) );
  COND2XL U2047 ( .A(n36), .B(n1306), .C(n1305), .D(n1658), .Z(n1022) );
  COND2XL U2048 ( .A(n36), .B(n1328), .C(n1327), .D(n1658), .Z(n1044) );
  COND2XL U2049 ( .A(n36), .B(n1307), .C(n1306), .D(n1658), .Z(n1023) );
  COND2XL U2050 ( .A(n36), .B(n1308), .C(n1307), .D(n1658), .Z(n1024) );
  COND2XL U2051 ( .A(n36), .B(n1326), .C(n1325), .D(n1658), .Z(n1042) );
  COND2XL U2052 ( .A(n36), .B(n1330), .C(n1329), .D(n1658), .Z(n1046) );
  CNR2IXL U2053 ( .B(n1746), .A(n1658), .Z(n1047) );
  COND2XL U2054 ( .A(n36), .B(n1329), .C(n1328), .D(n1658), .Z(n1045) );
  COND2XL U2055 ( .A(n36), .B(n1323), .C(n1322), .D(n1658), .Z(n1039) );
  COND2XL U2056 ( .A(n36), .B(n1309), .C(n1308), .D(n1658), .Z(n1025) );
  COND2XL U2057 ( .A(n36), .B(n1319), .C(n1318), .D(n1658), .Z(n1035) );
  CENX1 U2058 ( .A(n1734), .B(n1699), .Z(n1326) );
  CENX1 U2059 ( .A(n1735), .B(n155), .Z(n1309) );
  CANR1XL U2060 ( .A(n320), .B(n329), .C(n321), .Z(n319) );
  COND1XL U2061 ( .A(n298), .B(n311), .C(n299), .Z(n297) );
  COND2XL U2062 ( .A(n61), .B(n1569), .C(n1256), .D(n1617), .Z(n859) );
  COND2XL U2063 ( .A(n18), .B(n1362), .C(n1632), .D(n1361), .Z(n1076) );
  COND2XL U2064 ( .A(n18), .B(n1725), .C(n1391), .D(n1632), .Z(n864) );
  COND2XL U2065 ( .A(n18), .B(n1363), .C(n1631), .D(n1362), .Z(n1077) );
  COND2XL U2066 ( .A(n18), .B(n1388), .C(n1631), .D(n1387), .Z(n1102) );
  COND2XL U2067 ( .A(n18), .B(n1385), .C(n1631), .D(n1384), .Z(n1099) );
  COND2XL U2068 ( .A(n18), .B(n1383), .C(n1632), .D(n1382), .Z(n1097) );
  COND2XL U2069 ( .A(n18), .B(n1390), .C(n1632), .D(n1389), .Z(n1104) );
  COND2XL U2070 ( .A(n18), .B(n1389), .C(n1632), .D(n1388), .Z(n1103) );
  COND2XL U2071 ( .A(n18), .B(n1386), .C(n1632), .D(n1385), .Z(n1100) );
  COND2XL U2072 ( .A(n18), .B(n1384), .C(n1631), .D(n1383), .Z(n1098) );
  COND2XL U2073 ( .A(n18), .B(n1375), .C(n1631), .D(n1374), .Z(n1089) );
  COND2XL U2074 ( .A(n18), .B(n1365), .C(n1632), .D(n1364), .Z(n1079) );
  COND2XL U2075 ( .A(n18), .B(n1370), .C(n1631), .D(n1369), .Z(n1084) );
  COND2XL U2076 ( .A(n18), .B(n1379), .C(n1631), .D(n1378), .Z(n1093) );
  COND2XL U2077 ( .A(n18), .B(n1369), .C(n1632), .D(n1368), .Z(n1083) );
  COND2X1 U2078 ( .A(n18), .B(n1373), .C(n1632), .D(n1372), .Z(n1087) );
  CENX1 U2079 ( .A(n1736), .B(n151), .Z(n1313) );
  CENX1 U2080 ( .A(n1745), .B(n1736), .Z(n1330) );
  CND2XL U2081 ( .A(n653), .B(n672), .Z(n1687) );
  CND2X1 U2082 ( .A(n653), .B(n655), .Z(n1688) );
  CND2XL U2083 ( .A(n672), .B(n655), .Z(n1689) );
  COND2XL U2084 ( .A(n69), .B(n1218), .C(n1217), .D(n66), .Z(n938) );
  COND2XL U2085 ( .A(n69), .B(n1219), .C(n1218), .D(n66), .Z(n939) );
  COND2XL U2086 ( .A(n69), .B(n1221), .C(n1220), .D(n66), .Z(n941) );
  CNR2IXL U2087 ( .B(n1746), .A(n66), .Z(n955) );
  COND2XL U2088 ( .A(n69), .B(n1226), .C(n1225), .D(n66), .Z(n946) );
  COND2XL U2089 ( .A(n69), .B(n1227), .C(n1226), .D(n66), .Z(n947) );
  COND2XL U2090 ( .A(n69), .B(n1225), .C(n1224), .D(n66), .Z(n945) );
  COND2XL U2091 ( .A(n69), .B(n1232), .C(n1231), .D(n66), .Z(n952) );
  COND2XL U2092 ( .A(n69), .B(n1639), .C(n66), .D(n1235), .Z(n858) );
  COND2XL U2093 ( .A(n69), .B(n1224), .C(n1223), .D(n66), .Z(n944) );
  CIVX1 U2094 ( .A(n1725), .Z(n1719) );
  CIVX1 U2095 ( .A(n1725), .Z(n1724) );
  CIVX1 U2096 ( .A(n1725), .Z(n1721) );
  CIVX1 U2097 ( .A(n1742), .Z(n1740) );
  COND2XL U2098 ( .A(n36), .B(n1737), .C(n1331), .D(n1658), .Z(n862) );
  CND2IXL U2099 ( .B(n1746), .A(n1733), .Z(n1331) );
  CENX1 U2100 ( .A(n1733), .B(n156), .Z(n1308) );
  CENX1 U2101 ( .A(n1733), .B(n153), .Z(n1311) );
  COND2XL U2102 ( .A(n9), .B(n1565), .C(n6), .D(n1424), .Z(n865) );
  CND2X1 U2103 ( .A(n589), .B(n591), .Z(n1690) );
  CND2XL U2104 ( .A(n589), .B(n610), .Z(n1691) );
  CND2XL U2105 ( .A(n591), .B(n610), .Z(n1692) );
  CND3XL U2106 ( .A(n1690), .B(n1691), .C(n1692), .Z(n586) );
  CNR2X1 U2107 ( .A(n563), .B(n586), .Z(n239) );
  CEOX1 U2108 ( .A(a[6]), .B(n1736), .Z(n1455) );
  CIVX1 U2109 ( .A(n1737), .Z(n1736) );
  CEOXL U2110 ( .A(n360), .B(n190), .Z(product[7]) );
  CEOXL U2111 ( .A(n368), .B(n192), .Z(product[5]) );
  CND2XL U2112 ( .A(n489), .B(n491), .Z(n1693) );
  CND2XL U2113 ( .A(n489), .B(n514), .Z(n1694) );
  CND2X1 U2114 ( .A(n491), .B(n514), .Z(n1695) );
  CND3XL U2115 ( .A(n1693), .B(n1694), .C(n1695), .Z(n486) );
  CIVXL U2116 ( .A(n1725), .Z(n1722) );
  CIVXL U2117 ( .A(n1732), .Z(n1726) );
  CIVXL U2118 ( .A(n1732), .Z(n1728) );
  CIVXL U2119 ( .A(n1732), .Z(n1729) );
  CIVXL U2120 ( .A(n1732), .Z(n1730) );
  CIVXL U2121 ( .A(n1732), .Z(n1731) );
  CIVX2 U2122 ( .A(n21), .Z(n1732) );
  CIVXL U2123 ( .A(n1737), .Z(n1733) );
  CIVX2 U2124 ( .A(n374), .Z(n412) );
  CIVX2 U2125 ( .A(n336), .Z(n404) );
  CIVX2 U2126 ( .A(n333), .Z(n403) );
  CIVX2 U2127 ( .A(n322), .Z(n401) );
  CIVX2 U2128 ( .A(n295), .Z(n397) );
  CIVX2 U2129 ( .A(n223), .Z(n388) );
  CIVX2 U2130 ( .A(n218), .Z(n387) );
  CIVX2 U2131 ( .A(n383), .Z(n381) );
  CIVX2 U2132 ( .A(n380), .Z(n378) );
  CIVX2 U2133 ( .A(n372), .Z(n370) );
  CIVX2 U2134 ( .A(n364), .Z(n362) );
  CIVX2 U2135 ( .A(n356), .Z(n354) );
  CIVX2 U2136 ( .A(n352), .Z(n351) );
  CIVX2 U2137 ( .A(n350), .Z(n348) );
  CIVX2 U2138 ( .A(n345), .Z(n343) );
  CIVX2 U2139 ( .A(n328), .Z(n326) );
  CIVX2 U2140 ( .A(n327), .Z(n402) );
  CIVX2 U2141 ( .A(n318), .Z(n316) );
  CIVX2 U2142 ( .A(n306), .Z(n308) );
  CIVX2 U2143 ( .A(n305), .Z(n399) );
  CIVX2 U2144 ( .A(n290), .Z(n288) );
  CIVX2 U2145 ( .A(n285), .Z(n283) );
  CIVX2 U2146 ( .A(n273), .Z(n275) );
  CIVX2 U2147 ( .A(n272), .Z(n394) );
  CIVX2 U2148 ( .A(n250), .Z(n248) );
  CIVX2 U2149 ( .A(n1714), .Z(n1473) );
  CIVX2 U2150 ( .A(n1717), .Z(n1470) );
  CIVX2 U2151 ( .A(n113), .Z(n1468) );
endmodule


module calc_DW_mult_uns_19 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n89, n90, n92, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n108, n109, n110, n111, n113, n116, n117,
         n118, n120, n121, n122, n123, n124, n125, n126, n127, n128, n130,
         n132, n133, n134, n135, n139, n141, n142, n143, n144, n145, n146,
         n150, n152, n153, n154, n155, n157, n160, n161, n162, n163, n165,
         n167, n168, n170, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n184, n185, n186, n187, n188, n193, n194, n195, n196,
         n198, n200, n201, n203, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n220, n222, n223, n225,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n243, n245, n246, n247, n248, n251, n252,
         n253, n255, n257, n258, n261, n264, n265, n266, n267, n271, n274,
         n275, n276, n279, n280, n283, n284, n285, n287, n288, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n936, n961, n962, n963, \b[0] , n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070;
  assign product[0] = \b[0] ;
  assign \b[0]  = b[0];

  CEO3X2 U314 ( .A(n299), .B(n319), .C(n317), .Z(n295) );
  CEO3X2 U315 ( .A(n301), .B(n300), .C(n321), .Z(n296) );
  CEO3X2 U316 ( .A(n325), .B(n302), .C(n303), .Z(n297) );
  CEO3X2 U317 ( .A(n304), .B(n329), .C(n327), .Z(n298) );
  CEO3X2 U318 ( .A(n697), .B(n331), .C(n323), .Z(n299) );
  CEO3X2 U319 ( .A(n763), .B(n733), .C(n742), .Z(n300) );
  CEO3X2 U320 ( .A(n752), .B(n707), .C(n703), .Z(n301) );
  CEO3X2 U321 ( .A(n775), .B(n725), .C(n700), .Z(n302) );
  CEO3X2 U322 ( .A(n788), .B(n718), .C(n698), .Z(n303) );
  CFA1X1 U324 ( .A(n310), .B(n308), .CI(n335), .CO(n305), .S(n306) );
  CFA1X1 U325 ( .A(n339), .B(n337), .CI(n312), .CO(n307), .S(n308) );
  CFA1X1 U326 ( .A(n316), .B(n314), .CI(n341), .CO(n309), .S(n310) );
  CFA1X1 U327 ( .A(n320), .B(n318), .CI(n343), .CO(n311), .S(n312) );
  CFA1X1 U328 ( .A(n322), .B(n345), .CI(n347), .CO(n313), .S(n314) );
  CFA1X1 U329 ( .A(n328), .B(n324), .CI(n326), .CO(n315), .S(n316) );
  CFA1X1 U330 ( .A(n355), .B(n330), .CI(n349), .CO(n317), .S(n318) );
  CFA1X1 U331 ( .A(n332), .B(n353), .CI(n351), .CO(n319), .S(n320) );
  CFA1X1 U332 ( .A(n753), .B(n357), .CI(n699), .CO(n321), .S(n322) );
  CFA1X1 U333 ( .A(n776), .B(n734), .CI(n743), .CO(n323), .S(n324) );
  CFA1X1 U334 ( .A(n817), .B(n708), .CI(n726), .CO(n325), .S(n326) );
  CFA1X1 U335 ( .A(n764), .B(n704), .CI(n713), .CO(n327), .S(n328) );
  CFA1X1 U336 ( .A(n803), .B(n701), .CI(n719), .CO(n329), .S(n330) );
  CHA1X1 U337 ( .A(a[15]), .B(n789), .CO(n331), .S(n332) );
  CFA1X1 U338 ( .A(n338), .B(n336), .CI(n361), .CO(n333), .S(n334) );
  CFA1X1 U339 ( .A(n342), .B(n363), .CI(n340), .CO(n335), .S(n336) );
  CFA1X1 U340 ( .A(n367), .B(n365), .CI(n344), .CO(n337), .S(n338) );
  CFA1X1 U341 ( .A(n348), .B(n346), .CI(n369), .CO(n339), .S(n340) );
  CFA1X1 U342 ( .A(n354), .B(n371), .CI(n350), .CO(n341), .S(n342) );
  CFA1X1 U343 ( .A(n356), .B(n373), .CI(n352), .CO(n343), .S(n344) );
  CFA1X1 U344 ( .A(n375), .B(n381), .CI(n379), .CO(n345), .S(n346) );
  CFA1X1 U345 ( .A(n383), .B(n377), .CI(n358), .CO(n347), .S(n348) );
  CFA1X1 U346 ( .A(n765), .B(n702), .CI(n754), .CO(n349), .S(n350) );
  CFA1X1 U347 ( .A(n790), .B(n709), .CI(n744), .CO(n351), .S(n352) );
  CFA1X1 U348 ( .A(n818), .B(n714), .CI(n735), .CO(n353), .S(n354) );
  CFA1X1 U349 ( .A(n777), .B(n705), .CI(n727), .CO(n355), .S(n356) );
  CHA1X1 U350 ( .A(n804), .B(n720), .CO(n357), .S(n358) );
  CFA1X1 U351 ( .A(n364), .B(n362), .CI(n387), .CO(n359), .S(n360) );
  CFA1X1 U352 ( .A(n391), .B(n389), .CI(n366), .CO(n361), .S(n362) );
  CFA1X1 U353 ( .A(n393), .B(n368), .CI(n370), .CO(n363), .S(n364) );
  CFA1X1 U354 ( .A(n397), .B(n372), .CI(n395), .CO(n365), .S(n366) );
  CFA1X1 U355 ( .A(n382), .B(n374), .CI(n380), .CO(n367), .S(n368) );
  CFA1X1 U356 ( .A(n399), .B(n376), .CI(n378), .CO(n369), .S(n370) );
  CFA1X1 U357 ( .A(n403), .B(n405), .CI(n401), .CO(n371), .S(n372) );
  CFA1X1 U358 ( .A(n706), .B(n384), .CI(n407), .CO(n373), .S(n374) );
  CFA1X1 U359 ( .A(n778), .B(n755), .CI(n766), .CO(n375), .S(n376) );
  CFA1X1 U360 ( .A(n832), .B(n721), .CI(n745), .CO(n377), .S(n378) );
  CFA1X1 U361 ( .A(n805), .B(n715), .CI(n736), .CO(n379), .S(n380) );
  CFA1X1 U362 ( .A(n819), .B(n710), .CI(n728), .CO(n381), .S(n382) );
  CHA1X1 U363 ( .A(a[14]), .B(n791), .CO(n383), .S(n384) );
  CFA1X1 U364 ( .A(n390), .B(n388), .CI(n411), .CO(n385), .S(n386) );
  CFA1X1 U365 ( .A(n415), .B(n413), .CI(n392), .CO(n387), .S(n388) );
  CFA1X1 U366 ( .A(n417), .B(n394), .CI(n396), .CO(n389), .S(n390) );
  CFA1X1 U367 ( .A(n421), .B(n398), .CI(n419), .CO(n391), .S(n392) );
  CFA1X1 U368 ( .A(n404), .B(n400), .CI(n402), .CO(n393), .S(n394) );
  CFA1X1 U369 ( .A(n427), .B(n406), .CI(n423), .CO(n395), .S(n396) );
  CFA1X1 U370 ( .A(n408), .B(n429), .CI(n425), .CO(n397), .S(n398) );
  CFA1X1 U371 ( .A(n779), .B(n431), .CI(n711), .CO(n399), .S(n400) );
  CFA1X1 U372 ( .A(n792), .B(n729), .CI(n767), .CO(n401), .S(n402) );
  CFA1X1 U373 ( .A(n833), .B(n722), .CI(n756), .CO(n403), .S(n404) );
  CFA1X1 U374 ( .A(n820), .B(n716), .CI(n746), .CO(n405), .S(n406) );
  CHA1X1 U375 ( .A(n806), .B(n737), .CO(n407), .S(n408) );
  CFA1X1 U376 ( .A(n414), .B(n412), .CI(n435), .CO(n409), .S(n410) );
  CFA1X1 U377 ( .A(n439), .B(n437), .CI(n416), .CO(n411), .S(n412) );
  CFA1X1 U378 ( .A(n441), .B(n418), .CI(n420), .CO(n413), .S(n414) );
  CFA1X1 U379 ( .A(n445), .B(n422), .CI(n443), .CO(n415), .S(n416) );
  CFA1X1 U380 ( .A(n428), .B(n424), .CI(n426), .CO(n417), .S(n418) );
  CFA1X1 U381 ( .A(n447), .B(n430), .CI(n451), .CO(n419), .S(n420) );
  CFA1X1 U382 ( .A(n453), .B(n449), .CI(n432), .CO(n421), .S(n422) );
  CFA1X1 U383 ( .A(n846), .B(n717), .CI(n780), .CO(n423), .S(n424) );
  CFA1X1 U384 ( .A(n807), .B(n757), .CI(n768), .CO(n425), .S(n426) );
  CFA1X1 U385 ( .A(n793), .B(n738), .CI(n730), .CO(n427), .S(n428) );
  CFA1X1 U386 ( .A(n834), .B(n723), .CI(n747), .CO(n429), .S(n430) );
  CFA1X1 U388 ( .A(n438), .B(n436), .CI(n457), .CO(n433), .S(n434) );
  CFA1X1 U389 ( .A(n461), .B(n459), .CI(n440), .CO(n435), .S(n436) );
  CFA1X1 U390 ( .A(n463), .B(n442), .CI(n444), .CO(n437), .S(n438) );
  CFA1X1 U391 ( .A(n450), .B(n446), .CI(n465), .CO(n439), .S(n440) );
  CFA1X1 U392 ( .A(n452), .B(n467), .CI(n448), .CO(n441), .S(n442) );
  CFA1X1 U393 ( .A(n469), .B(n473), .CI(n471), .CO(n443), .S(n444) );
  CFA1X1 U394 ( .A(n724), .B(n454), .CI(n475), .CO(n445), .S(n446) );
  CFA1X1 U395 ( .A(n847), .B(n794), .CI(n781), .CO(n447), .S(n448) );
  CFA1X1 U396 ( .A(n822), .B(n758), .CI(n769), .CO(n449), .S(n450) );
  CFA1X1 U397 ( .A(n808), .B(n731), .CI(n748), .CO(n451), .S(n452) );
  CHA1X1 U398 ( .A(n835), .B(n739), .CO(n453), .S(n454) );
  CFA1X1 U399 ( .A(n460), .B(n458), .CI(n479), .CO(n455), .S(n456) );
  CFA1X1 U400 ( .A(n464), .B(n481), .CI(n462), .CO(n457), .S(n458) );
  CFA1X1 U401 ( .A(n485), .B(n483), .CI(n466), .CO(n459), .S(n460) );
  CFA1X1 U402 ( .A(n472), .B(n487), .CI(n468), .CO(n461), .S(n462) );
  CFA1X1 U403 ( .A(n489), .B(n470), .CI(n474), .CO(n463), .S(n464) );
  CFA1X1 U404 ( .A(n476), .B(n493), .CI(n491), .CO(n465), .S(n466) );
  CFA1X1 U405 ( .A(n809), .B(n495), .CI(n732), .CO(n467), .S(n468) );
  CFA1X1 U406 ( .A(n859), .B(n782), .CI(n795), .CO(n469), .S(n470) );
  CFA1X1 U407 ( .A(n848), .B(n759), .CI(n770), .CO(n471), .S(n472) );
  CFA1X1 U408 ( .A(n823), .B(n740), .CI(n749), .CO(n473), .S(n474) );
  CFA1X1 U410 ( .A(n482), .B(n480), .CI(n499), .CO(n477), .S(n478) );
  CFA1X1 U411 ( .A(n486), .B(n501), .CI(n484), .CO(n479), .S(n480) );
  CFA1X1 U412 ( .A(n505), .B(n503), .CI(n488), .CO(n481), .S(n482) );
  CFA1X1 U413 ( .A(n494), .B(n507), .CI(n490), .CO(n483), .S(n484) );
  CFA1X1 U414 ( .A(n509), .B(n492), .CI(n513), .CO(n485), .S(n486) );
  CFA1X1 U415 ( .A(n515), .B(n511), .CI(n496), .CO(n487), .S(n488) );
  CFA1X1 U416 ( .A(n824), .B(n741), .CI(n810), .CO(n489), .S(n490) );
  CFA1X1 U417 ( .A(n849), .B(n783), .CI(n796), .CO(n491), .S(n492) );
  CFA1X1 U418 ( .A(n860), .B(n771), .CI(n760), .CO(n493), .S(n494) );
  CHA1X1 U419 ( .A(n837), .B(n750), .CO(n495), .S(n496) );
  CFA1X1 U420 ( .A(n502), .B(n500), .CI(n519), .CO(n497), .S(n498) );
  CFA1X1 U421 ( .A(n506), .B(n521), .CI(n504), .CO(n499), .S(n500) );
  CFA1X1 U422 ( .A(n508), .B(n523), .CI(n525), .CO(n501), .S(n502) );
  CFA1X1 U423 ( .A(n514), .B(n510), .CI(n512), .CO(n503), .S(n504) );
  CFA1X1 U424 ( .A(n529), .B(n527), .CI(n531), .CO(n505), .S(n506) );
  CFA1X1 U425 ( .A(n751), .B(n516), .CI(n533), .CO(n507), .S(n508) );
  CFA1X1 U426 ( .A(n838), .B(n811), .CI(n825), .CO(n509), .S(n510) );
  CFA1X1 U427 ( .A(n871), .B(n784), .CI(n797), .CO(n511), .S(n512) );
  CFA1X1 U428 ( .A(n850), .B(n761), .CI(n772), .CO(n513), .S(n514) );
  CFA1X1 U430 ( .A(n522), .B(n520), .CI(n537), .CO(n517), .S(n518) );
  CFA1X1 U431 ( .A(n541), .B(n539), .CI(n524), .CO(n519), .S(n520) );
  CFA1X1 U432 ( .A(n528), .B(n526), .CI(n543), .CO(n521), .S(n522) );
  CFA1X1 U433 ( .A(n545), .B(n532), .CI(n530), .CO(n523), .S(n524) );
  CFA1X1 U434 ( .A(n534), .B(n549), .CI(n547), .CO(n525), .S(n526) );
  CFA1X1 U435 ( .A(n872), .B(n551), .CI(n762), .CO(n527), .S(n528) );
  CFA1X1 U436 ( .A(n851), .B(n812), .CI(n826), .CO(n529), .S(n530) );
  CFA1X1 U437 ( .A(n839), .B(n798), .CI(n785), .CO(n531), .S(n532) );
  CHA1X1 U438 ( .A(n862), .B(n773), .CO(n533), .S(n534) );
  CFA1X1 U439 ( .A(n540), .B(n538), .CI(n555), .CO(n535), .S(n536) );
  CFA1X1 U440 ( .A(n544), .B(n557), .CI(n542), .CO(n537), .S(n538) );
  CFA1X1 U441 ( .A(n546), .B(n559), .CI(n561), .CO(n539), .S(n540) );
  CFA1X1 U442 ( .A(n565), .B(n550), .CI(n548), .CO(n541), .S(n542) );
  CFA1X1 U443 ( .A(n567), .B(n563), .CI(n552), .CO(n543), .S(n544) );
  CFA1X1 U444 ( .A(n873), .B(n774), .CI(n840), .CO(n545), .S(n546) );
  CFA1X1 U445 ( .A(n852), .B(n813), .CI(n827), .CO(n547), .S(n548) );
  CFA1X1 U446 ( .A(n863), .B(n786), .CI(n799), .CO(n549), .S(n550) );
  CFA1X1 U448 ( .A(n558), .B(n556), .CI(n571), .CO(n553), .S(n554) );
  CFA1X1 U449 ( .A(n562), .B(n573), .CI(n560), .CO(n555), .S(n556) );
  CFA1X1 U450 ( .A(n564), .B(n575), .CI(n577), .CO(n557), .S(n558) );
  CFA1X1 U451 ( .A(n579), .B(n566), .CI(n581), .CO(n559), .S(n560) );
  CFA1X1 U452 ( .A(n787), .B(n568), .CI(n583), .CO(n561), .S(n562) );
  CFA1X1 U453 ( .A(n874), .B(n841), .CI(n853), .CO(n563), .S(n564) );
  CFA1X1 U454 ( .A(n864), .B(n828), .CI(n814), .CO(n565), .S(n566) );
  CHA1X1 U455 ( .A(n883), .B(n800), .CO(n567), .S(n568) );
  CFA1X1 U456 ( .A(n574), .B(n572), .CI(n587), .CO(n569), .S(n570) );
  CFA1X1 U457 ( .A(n591), .B(n589), .CI(n576), .CO(n571), .S(n572) );
  CFA1X1 U458 ( .A(n582), .B(n578), .CI(n580), .CO(n573), .S(n574) );
  CFA1X1 U459 ( .A(n584), .B(n593), .CI(n595), .CO(n575), .S(n576) );
  CFA1X1 U460 ( .A(n854), .B(n597), .CI(n801), .CO(n577), .S(n578) );
  CFA1X1 U461 ( .A(n865), .B(n842), .CI(n892), .CO(n579), .S(n580) );
  CFA1X1 U462 ( .A(n875), .B(n815), .CI(n829), .CO(n581), .S(n582) );
  CFA1X1 U464 ( .A(n590), .B(n588), .CI(n601), .CO(n585), .S(n586) );
  CFA1X1 U465 ( .A(n605), .B(n603), .CI(n592), .CO(n587), .S(n588) );
  CFA1X1 U466 ( .A(n607), .B(n594), .CI(n596), .CO(n589), .S(n590) );
  CFA1X1 U467 ( .A(n611), .B(n609), .CI(n598), .CO(n591), .S(n592) );
  CFA1X1 U468 ( .A(n866), .B(n816), .CI(n893), .CO(n593), .S(n594) );
  CFA1X1 U469 ( .A(n876), .B(n855), .CI(n843), .CO(n595), .S(n596) );
  CHA1X1 U470 ( .A(n885), .B(n830), .CO(n597), .S(n598) );
  CFA1X1 U471 ( .A(n604), .B(n602), .CI(n615), .CO(n599), .S(n600) );
  CFA1X1 U472 ( .A(n608), .B(n617), .CI(n606), .CO(n601), .S(n602) );
  CFA1X1 U473 ( .A(n621), .B(n610), .CI(n619), .CO(n603), .S(n604) );
  CFA1X1 U474 ( .A(n831), .B(n612), .CI(n623), .CO(n605), .S(n606) );
  CFA1X1 U475 ( .A(n901), .B(n867), .CI(n894), .CO(n607), .S(n608) );
  CFA1X1 U476 ( .A(n877), .B(n844), .CI(n856), .CO(n609), .S(n610) );
  CFA1X1 U478 ( .A(n618), .B(n616), .CI(n627), .CO(n613), .S(n614) );
  CFA1X1 U479 ( .A(n622), .B(n629), .CI(n620), .CO(n615), .S(n616) );
  CFA1X1 U480 ( .A(n624), .B(n631), .CI(n633), .CO(n617), .S(n618) );
  CFA1X1 U481 ( .A(n895), .B(n635), .CI(n845), .CO(n619), .S(n620) );
  CFA1X1 U482 ( .A(n902), .B(n868), .CI(n878), .CO(n621), .S(n622) );
  CHA1X1 U483 ( .A(n887), .B(n857), .CO(n623), .S(n624) );
  CFA1X1 U484 ( .A(n630), .B(n628), .CI(n639), .CO(n625), .S(n626) );
  CFA1X1 U485 ( .A(n634), .B(n641), .CI(n632), .CO(n627), .S(n628) );
  CFA1X1 U486 ( .A(n645), .B(n643), .CI(n636), .CO(n629), .S(n630) );
  CFA1X1 U487 ( .A(n888), .B(n858), .CI(n879), .CO(n631), .S(n632) );
  CFA1X1 U488 ( .A(n903), .B(n869), .CI(n909), .CO(n633), .S(n634) );
  CFA1X1 U490 ( .A(n642), .B(n640), .CI(n649), .CO(n637), .S(n638) );
  CFA1X1 U491 ( .A(n653), .B(n644), .CI(n651), .CO(n639), .S(n640) );
  CFA1X1 U492 ( .A(n870), .B(n646), .CI(n655), .CO(n641), .S(n642) );
  CFA1X1 U493 ( .A(n889), .B(n910), .CI(n897), .CO(n643), .S(n644) );
  CHA1X1 U494 ( .A(n904), .B(n880), .CO(n645), .S(n646) );
  CFA1X1 U495 ( .A(n652), .B(n650), .CI(n659), .CO(n647), .S(n648) );
  CFA1X1 U496 ( .A(n656), .B(n654), .CI(n661), .CO(n649), .S(n650) );
  CFA1X1 U497 ( .A(n916), .B(n663), .CI(n881), .CO(n651), .S(n652) );
  CFA1X1 U498 ( .A(n898), .B(n890), .CI(n911), .CO(n653), .S(n654) );
  CFA1X1 U500 ( .A(n662), .B(n660), .CI(n667), .CO(n657), .S(n658) );
  CFA1X1 U501 ( .A(n671), .B(n669), .CI(n664), .CO(n659), .S(n660) );
  CFA1X1 U502 ( .A(n917), .B(n891), .CI(n912), .CO(n661), .S(n662) );
  CHA1X1 U503 ( .A(n906), .B(n899), .CO(n663), .S(n664) );
  CFA1X1 U504 ( .A(n675), .B(n668), .CI(n670), .CO(n665), .S(n666) );
  CFA1X1 U505 ( .A(n900), .B(n672), .CI(n677), .CO(n667), .S(n668) );
  CFA1X1 U506 ( .A(n913), .B(n907), .CI(n922), .CO(n669), .S(n670) );
  CHA1X1 U507 ( .A(a[5]), .B(n918), .CO(n671), .S(n672) );
  CFA1X1 U508 ( .A(n678), .B(n676), .CI(n681), .CO(n673), .S(n674) );
  CFA1X1 U509 ( .A(n923), .B(n683), .CI(n908), .CO(n675), .S(n676) );
  CHA1X1 U510 ( .A(n919), .B(n914), .CO(n677), .S(n678) );
  CFA1X1 U511 ( .A(n687), .B(n682), .CI(n684), .CO(n679), .S(n680) );
  CFA1X1 U512 ( .A(n920), .B(n915), .CI(n927), .CO(n681), .S(n682) );
  CFA1X1 U514 ( .A(n921), .B(n688), .CI(n691), .CO(n685), .S(n686) );
  CHA1X1 U515 ( .A(n925), .B(n928), .CO(n687), .S(n688) );
  CFA1X1 U516 ( .A(n931), .B(n692), .CI(n926), .CO(n689), .S(n690) );
  CHA1X1 U518 ( .A(n932), .B(n930), .CO(n693), .S(n694) );
  COND1X1 U808 ( .A(n122), .B(n116), .C(n117), .Z(n111) );
  CIVX2 U809 ( .A(b[21]), .Z(n21) );
  CNR2X1 U810 ( .A(n1058), .B(n961), .Z(n843) );
  CNR2X1 U811 ( .A(n1067), .B(n15), .Z(n822) );
  CIVX2 U812 ( .A(b[11]), .Z(n1070) );
  CIVX2 U813 ( .A(b[12]), .Z(n963) );
  CANR1XL U814 ( .A(n238), .B(n230), .C(n231), .Z(n229) );
  COND1XL U815 ( .A(n162), .B(n174), .C(n163), .Z(n161) );
  CANR1XL U816 ( .A(n170), .B(n1042), .C(n165), .Z(n163) );
  CIVX2 U817 ( .A(b[8]), .Z(n1065) );
  CIVX2 U818 ( .A(b[3]), .Z(n1060) );
  CIVX2 U819 ( .A(b[5]), .Z(n1062) );
  CIVX2 U820 ( .A(b[6]), .Z(n1063) );
  CIVX2 U821 ( .A(b[10]), .Z(n1068) );
  CIVX2 U822 ( .A(b[9]), .Z(n1067) );
  CIVX1 U823 ( .A(b[9]), .Z(n1066) );
  CIVX2 U824 ( .A(b[4]), .Z(n1061) );
  CIVX2 U825 ( .A(b[7]), .Z(n1064) );
  CAN2X1 U826 ( .A(n1038), .B(n261), .Z(product[2]) );
  CIVXL U827 ( .A(n161), .Z(n160) );
  CIVXL U828 ( .A(b[25]), .Z(n25) );
  CNR2XL U829 ( .A(n1057), .B(n1063), .Z(n920) );
  CIVX3 U830 ( .A(b[13]), .Z(n962) );
  COR2X1 U831 ( .A(n658), .B(n665), .Z(n1047) );
  CNR2XL U832 ( .A(n1058), .B(n1069), .Z(n879) );
  CNR2XL U833 ( .A(n1059), .B(n1064), .Z(n913) );
  CIVX2 U834 ( .A(b[16]), .Z(n16) );
  CND2XL U835 ( .A(n1039), .B(n94), .Z(n60) );
  CANR1X1 U836 ( .A(n208), .B(n216), .C(n209), .Z(n207) );
  CNR2XL U837 ( .A(n232), .B(n235), .Z(n230) );
  CNR2XL U838 ( .A(n1064), .B(n1065), .Z(n901) );
  CNR2XL U839 ( .A(n1063), .B(n1064), .Z(n909) );
  CNR2XL U840 ( .A(n963), .B(n15), .Z(n819) );
  CNR2XL U841 ( .A(n1061), .B(n1063), .Z(n917) );
  CNR2XL U842 ( .A(n1060), .B(n1064), .Z(n912) );
  CNR2XL U843 ( .A(n1054), .B(n1068), .Z(n891) );
  CNR2XL U844 ( .A(n1057), .B(n1065), .Z(n907) );
  CNR2XL U845 ( .A(n1062), .B(n963), .Z(n865) );
  CNR2XL U846 ( .A(n1055), .B(n1062), .Z(n926) );
  CIVX2 U847 ( .A(b[14]), .Z(n961) );
  CIVXL U848 ( .A(b[26]), .Z(n26) );
  CENX1 U849 ( .A(n95), .B(n60), .Z(product[30]) );
  CNR2X1 U850 ( .A(n498), .B(n517), .Z(n154) );
  COR2X1 U851 ( .A(n536), .B(n553), .Z(n1044) );
  CND2XL U852 ( .A(n287), .B(n248), .Z(n84) );
  CANR1XL U853 ( .A(n258), .B(n1053), .C(n255), .Z(n253) );
  CNR2XL U854 ( .A(n1063), .B(n962), .Z(n852) );
  CNR2X1 U855 ( .A(n1070), .B(n16), .Z(n805) );
  CNR2XL U856 ( .A(n1061), .B(n963), .Z(n866) );
  CNR2XL U857 ( .A(n1063), .B(n1068), .Z(n885) );
  CNR2XL U858 ( .A(n1062), .B(n1063), .Z(n916) );
  CNR2XL U859 ( .A(n1062), .B(n961), .Z(n840) );
  CNR2X1 U860 ( .A(n1060), .B(n23), .Z(n729) );
  CNR2X1 U861 ( .A(n1054), .B(n1065), .Z(n908) );
  CNR2XL U862 ( .A(n1061), .B(n962), .Z(n854) );
  CNR2X1 U863 ( .A(n1065), .B(n18), .Z(n779) );
  CNR2X1 U864 ( .A(n1066), .B(n18), .Z(n778) );
  CEO3X1 U865 ( .A(n309), .B(n292), .C(n307), .Z(n291) );
  CEO3X1 U866 ( .A(n311), .B(n294), .C(n293), .Z(n292) );
  CEO3X1 U867 ( .A(n298), .B(n297), .C(n315), .Z(n294) );
  CEO3X1 U868 ( .A(n296), .B(n313), .C(n295), .Z(n293) );
  CIVX2 U869 ( .A(b[15]), .Z(n15) );
  CIVX2 U870 ( .A(b[17]), .Z(n17) );
  CNR2X1 U871 ( .A(n1057), .B(n1061), .Z(n929) );
  CANR1X1 U872 ( .A(n1039), .B(n95), .C(n92), .Z(n90) );
  COND1X1 U873 ( .A(n124), .B(n96), .C(n97), .Z(n95) );
  CNR2XL U874 ( .A(n116), .B(n121), .Z(n110) );
  CEOXL U875 ( .A(n62), .B(n109), .Z(product[28]) );
  CND2XL U876 ( .A(n265), .B(n108), .Z(n62) );
  CEOXL U877 ( .A(n61), .B(n102), .Z(product[29]) );
  CND2XL U878 ( .A(n267), .B(n122), .Z(n64) );
  CNR2IXL U879 ( .B(n110), .A(n105), .Z(n103) );
  CANR1X1 U880 ( .A(n161), .B(n125), .C(n126), .Z(n124) );
  CNR2XL U881 ( .A(n127), .B(n143), .Z(n125) );
  CND2XL U882 ( .A(n1043), .B(n1040), .Z(n127) );
  CND2XL U883 ( .A(n274), .B(n178), .Z(n71) );
  CND2XL U884 ( .A(n1040), .B(n141), .Z(n66) );
  CND2XL U885 ( .A(n1042), .B(n1044), .Z(n162) );
  CEOXL U886 ( .A(n69), .B(n168), .Z(product[21]) );
  CND2XL U887 ( .A(n1042), .B(n167), .Z(n69) );
  CEOXL U888 ( .A(n68), .B(n160), .Z(product[22]) );
  CND2XL U889 ( .A(n271), .B(n155), .Z(n68) );
  CND2XL U890 ( .A(n276), .B(n188), .Z(n73) );
  CND2XL U891 ( .A(n1041), .B(n152), .Z(n67) );
  CND2XL U892 ( .A(n1043), .B(n132), .Z(n65) );
  CND2XL U893 ( .A(n145), .B(n1040), .Z(n134) );
  CND2XL U894 ( .A(n1044), .B(n172), .Z(n70) );
  CND2XL U895 ( .A(n275), .B(n185), .Z(n72) );
  CND2XL U896 ( .A(n386), .B(n409), .Z(n117) );
  CND2XL U897 ( .A(n334), .B(n359), .Z(n101) );
  CANR1X1 U898 ( .A(n157), .B(n1041), .C(n150), .Z(n144) );
  CIVX1 U899 ( .A(n152), .Z(n150) );
  CNR2XL U900 ( .A(n210), .B(n213), .Z(n208) );
  CND2XL U901 ( .A(n1048), .B(n222), .Z(n78) );
  CND2XL U902 ( .A(n280), .B(n214), .Z(n77) );
  CND2XL U903 ( .A(n1045), .B(n200), .Z(n74) );
  CND2XL U904 ( .A(n570), .B(n585), .Z(n185) );
  CND2XL U905 ( .A(n1047), .B(n227), .Z(n79) );
  CND2XL U906 ( .A(n1046), .B(n205), .Z(n75) );
  CND2XL U907 ( .A(n666), .B(n673), .Z(n233) );
  CND2XL U908 ( .A(n626), .B(n637), .Z(n211) );
  CEOXL U909 ( .A(n1049), .B(n84), .Z(product[6]) );
  CND2XL U910 ( .A(n1050), .B(n245), .Z(n83) );
  CND2XL U911 ( .A(n283), .B(n233), .Z(n80) );
  CND2XL U912 ( .A(n284), .B(n236), .Z(n81) );
  CEOXL U913 ( .A(n59), .B(n90), .Z(product[31]) );
  CND2XL U914 ( .A(n680), .B(n685), .Z(n240) );
  CND2XL U915 ( .A(n690), .B(n693), .Z(n248) );
  CND2XL U916 ( .A(n288), .B(n252), .Z(n85) );
  CEOXL U917 ( .A(n253), .B(n85), .Z(product[5]) );
  CND2XL U918 ( .A(n1053), .B(n257), .Z(n86) );
  CNR2XL U919 ( .A(n1054), .B(n961), .Z(n845) );
  CNR2XL U920 ( .A(n1057), .B(n15), .Z(n830) );
  CNR2XL U921 ( .A(n1055), .B(n1064), .Z(n915) );
  CNR2XL U922 ( .A(n1060), .B(n1061), .Z(n927) );
  CNR2XL U923 ( .A(n1055), .B(n1063), .Z(n921) );
  CNR2XL U924 ( .A(n1058), .B(n962), .Z(n856) );
  CNR2XL U925 ( .A(n1061), .B(n1069), .Z(n877) );
  CNR2XL U926 ( .A(n1057), .B(n961), .Z(n844) );
  CNR2XL U927 ( .A(n1055), .B(n16), .Z(n816) );
  CNR2XL U928 ( .A(n1064), .B(n20), .Z(n755) );
  CNR2XL U929 ( .A(n1060), .B(n15), .Z(n828) );
  CNR2XL U930 ( .A(n1059), .B(n16), .Z(n814) );
  CNR2XL U931 ( .A(n1061), .B(n26), .Z(n707) );
  CNR2XL U932 ( .A(n1060), .B(n21), .Z(n748) );
  CNR2XL U933 ( .A(n1067), .B(n17), .Z(n792) );
  CNR2XL U934 ( .A(n1060), .B(n24), .Z(n721) );
  CNR2XL U935 ( .A(n1062), .B(n25), .Z(n712) );
  CNR2XL U936 ( .A(n1060), .B(n27), .Z(n703) );
  CNR2XL U937 ( .A(n1055), .B(n1057), .Z(n936) );
  CNR2XL U938 ( .A(n1054), .B(n1069), .Z(n881) );
  CNR2XL U939 ( .A(n1058), .B(n963), .Z(n868) );
  CNR2XL U940 ( .A(n1060), .B(n1069), .Z(n878) );
  CNR2XL U941 ( .A(n1060), .B(n963), .Z(n867) );
  CNR2XL U942 ( .A(n1054), .B(n21), .Z(n751) );
  CNR2XL U943 ( .A(n1055), .B(n19), .Z(n774) );
  CNR2XL U944 ( .A(n1060), .B(n20), .Z(n759) );
  CNR2XL U945 ( .A(n1061), .B(n19), .Z(n770) );
  CNR2XL U946 ( .A(n1055), .B(n20), .Z(n762) );
  CNR2XL U947 ( .A(n1057), .B(n963), .Z(n869) );
  CNR2XL U948 ( .A(n1060), .B(n22), .Z(n738) );
  CNR2XL U949 ( .A(n963), .B(n961), .Z(n833) );
  CNR2XL U950 ( .A(n1058), .B(n15), .Z(n829) );
  CNR2XL U951 ( .A(n1057), .B(n16), .Z(n815) );
  CNR2XL U952 ( .A(n1063), .B(n1069), .Z(n875) );
  CNR2XL U953 ( .A(n1068), .B(n18), .Z(n777) );
  CNR2XL U954 ( .A(n1062), .B(n23), .Z(n727) );
  CNR2XL U955 ( .A(n1057), .B(n27), .Z(n705) );
  CNR2XL U956 ( .A(n1060), .B(n25), .Z(n714) );
  CNR2XL U957 ( .A(n1061), .B(n20), .Z(n758) );
  CNR2XL U958 ( .A(n1066), .B(n20), .Z(n753) );
  CNR2XL U959 ( .A(n1068), .B(n19), .Z(n764) );
  CNR2XL U960 ( .A(n1058), .B(n27), .Z(n704) );
  CNR2XL U961 ( .A(n1061), .B(n25), .Z(n713) );
  CNR2XL U962 ( .A(n1060), .B(n16), .Z(n813) );
  CNR2XL U963 ( .A(n1054), .B(n18), .Z(n787) );
  CNR2XL U964 ( .A(n1065), .B(n963), .Z(n862) );
  CNR2XL U965 ( .A(n1057), .B(n962), .Z(n857) );
  CNR2XL U966 ( .A(n1061), .B(n1068), .Z(n887) );
  CNR2XL U967 ( .A(n1068), .B(n16), .Z(n806) );
  CNR2XL U968 ( .A(n1061), .B(n22), .Z(n737) );
  CNR2XL U969 ( .A(n1061), .B(n16), .Z(n812) );
  CNR2XL U970 ( .A(n1061), .B(n17), .Z(n797) );
  CNR2XL U971 ( .A(n1060), .B(n962), .Z(n855) );
  CNR2XL U972 ( .A(n1054), .B(n962), .Z(n858) );
  CNR2XL U973 ( .A(n1060), .B(n961), .Z(n842) );
  CNR2XL U974 ( .A(n1066), .B(n19), .Z(n765) );
  CNR2XL U975 ( .A(n1054), .B(n15), .Z(n831) );
  CNR2XL U976 ( .A(n1069), .B(n17), .Z(n790) );
  CNR2XL U977 ( .A(n1063), .B(n23), .Z(n726) );
  CNR2XL U978 ( .A(n1057), .B(n1067), .Z(n899) );
  CNR2XL U979 ( .A(n1061), .B(n24), .Z(n720) );
  CNR2XL U980 ( .A(n963), .B(n16), .Z(n804) );
  CNR2XL U981 ( .A(n1068), .B(n20), .Z(n752) );
  CNR2XL U982 ( .A(n963), .B(n18), .Z(n775) );
  CNR2XL U983 ( .A(n1054), .B(n963), .Z(n870) );
  COR2XL U984 ( .A(n1055), .B(n1058), .Z(n1052) );
  CNR2XL U985 ( .A(n1058), .B(n1068), .Z(n889) );
  CNR2XL U986 ( .A(n1062), .B(n1064), .Z(n910) );
  CNR2XL U987 ( .A(n1060), .B(n1062), .Z(n923) );
  CNR2XL U988 ( .A(n1055), .B(n17), .Z(n801) );
  CNR2XL U989 ( .A(n1061), .B(n18), .Z(n783) );
  CNR2XL U990 ( .A(n1061), .B(n21), .Z(n747) );
  CNR2XL U991 ( .A(n1054), .B(n24), .Z(n724) );
  CNR2XL U992 ( .A(n1070), .B(n18), .Z(n776) );
  CNR2XL U993 ( .A(n1059), .B(n1061), .Z(n928) );
  CNR2XL U994 ( .A(n1057), .B(n1062), .Z(n925) );
  CNR2XL U995 ( .A(n1059), .B(n1060), .Z(n931) );
  CNR2XL U996 ( .A(n1067), .B(n21), .Z(n742) );
  CNR2XL U997 ( .A(n1055), .B(n1061), .Z(n930) );
  CNR2XL U998 ( .A(n1057), .B(n1060), .Z(n932) );
  CEOXL U999 ( .A(n261), .B(n1052), .Z(product[3]) );
  CIVX1 U1000 ( .A(b[18]), .Z(n18) );
  CNR2XL U1001 ( .A(n1059), .B(n1062), .Z(n924) );
  CIVX1 U1002 ( .A(b[19]), .Z(n19) );
  CIVX1 U1003 ( .A(b[20]), .Z(n20) );
  CND2XL U1004 ( .A(n936), .B(a[1]), .Z(n261) );
  CIVXL U1005 ( .A(b[24]), .Z(n24) );
  CNR2XL U1006 ( .A(n963), .B(n17), .Z(n789) );
  CNR2XL U1007 ( .A(n1067), .B(n1068), .Z(n882) );
  COR2XL U1008 ( .A(n936), .B(a[1]), .Z(n1038) );
  CND2X1 U1009 ( .A(n98), .B(n110), .Z(n96) );
  CANR1XL U1010 ( .A(n111), .B(n98), .C(n99), .Z(n97) );
  CND2X1 U1011 ( .A(n266), .B(n117), .Z(n63) );
  CANR1XL U1012 ( .A(n267), .B(n123), .C(n120), .Z(n118) );
  CENX1 U1013 ( .A(n123), .B(n64), .Z(product[26]) );
  COND1XL U1014 ( .A(n108), .B(n100), .C(n101), .Z(n99) );
  COND1XL U1015 ( .A(n105), .B(n113), .C(n108), .Z(n104) );
  CANR1XL U1016 ( .A(n110), .B(n123), .C(n111), .Z(n109) );
  CND2X1 U1017 ( .A(n264), .B(n101), .Z(n61) );
  CANR1XL U1018 ( .A(n103), .B(n123), .C(n104), .Z(n102) );
  CND2X1 U1019 ( .A(n275), .B(n276), .Z(n180) );
  CNR2X1 U1020 ( .A(n360), .B(n385), .Z(n105) );
  CENX1 U1021 ( .A(n142), .B(n66), .Z(product[24]) );
  COND1XL U1022 ( .A(n144), .B(n127), .C(n128), .Z(n126) );
  CNR2X1 U1023 ( .A(n386), .B(n409), .Z(n116) );
  CANR1XL U1024 ( .A(n194), .B(n175), .C(n176), .Z(n174) );
  CNR2X1 U1025 ( .A(n180), .B(n177), .Z(n175) );
  COND1XL U1026 ( .A(n177), .B(n181), .C(n178), .Z(n176) );
  CANR1XL U1027 ( .A(n1040), .B(n146), .C(n139), .Z(n135) );
  CNR2X1 U1028 ( .A(n410), .B(n433), .Z(n121) );
  CNR2X1 U1029 ( .A(n334), .B(n359), .Z(n100) );
  CANR1XL U1030 ( .A(n139), .B(n1043), .C(n130), .Z(n128) );
  CENX1 U1031 ( .A(n179), .B(n71), .Z(product[19]) );
  CENX1 U1032 ( .A(n153), .B(n67), .Z(product[23]) );
  COND1XL U1033 ( .A(n154), .B(n160), .C(n155), .Z(n153) );
  CENX1 U1034 ( .A(n133), .B(n65), .Z(product[25]) );
  COND1XL U1035 ( .A(n134), .B(n160), .C(n135), .Z(n133) );
  CENX1 U1036 ( .A(n186), .B(n72), .Z(product[18]) );
  COND1XL U1037 ( .A(n187), .B(n193), .C(n188), .Z(n186) );
  CENX1 U1038 ( .A(n173), .B(n70), .Z(product[20]) );
  CANR1XL U1039 ( .A(n1044), .B(n173), .C(n170), .Z(n168) );
  CEOX1 U1040 ( .A(n73), .B(n193), .Z(product[17]) );
  CND2X1 U1041 ( .A(n410), .B(n433), .Z(n122) );
  CND2X1 U1042 ( .A(n1041), .B(n271), .Z(n143) );
  CND2X1 U1043 ( .A(n360), .B(n385), .Z(n108) );
  CND2X1 U1044 ( .A(n306), .B(n333), .Z(n94) );
  COR2X1 U1045 ( .A(n306), .B(n333), .Z(n1039) );
  COND1XL U1046 ( .A(n229), .B(n217), .C(n218), .Z(n216) );
  CND2X1 U1047 ( .A(n1048), .B(n1047), .Z(n217) );
  CANR1XL U1048 ( .A(n225), .B(n1048), .C(n220), .Z(n218) );
  CNR2X1 U1049 ( .A(n554), .B(n569), .Z(n177) );
  COND1XL U1050 ( .A(n214), .B(n210), .C(n211), .Z(n209) );
  COND1X1 U1051 ( .A(n195), .B(n207), .C(n196), .Z(n194) );
  CND2X1 U1052 ( .A(n1045), .B(n1046), .Z(n195) );
  CANR1XL U1053 ( .A(n203), .B(n1045), .C(n198), .Z(n196) );
  COR2X1 U1054 ( .A(n456), .B(n477), .Z(n1040) );
  CENX1 U1055 ( .A(n228), .B(n79), .Z(product[11]) );
  CENX1 U1056 ( .A(n212), .B(n76), .Z(product[14]) );
  CND2X1 U1057 ( .A(n279), .B(n211), .Z(n76) );
  COND1XL U1058 ( .A(n213), .B(n215), .C(n214), .Z(n212) );
  CENX1 U1059 ( .A(n206), .B(n75), .Z(product[15]) );
  CNR2X1 U1060 ( .A(n570), .B(n585), .Z(n184) );
  CEOX1 U1061 ( .A(n78), .B(n223), .Z(product[12]) );
  CANR1XL U1062 ( .A(n1047), .B(n228), .C(n225), .Z(n223) );
  CEOX1 U1063 ( .A(n77), .B(n215), .Z(product[13]) );
  CEOX1 U1064 ( .A(n74), .B(n201), .Z(product[16]) );
  CANR1XL U1065 ( .A(n1046), .B(n206), .C(n203), .Z(n201) );
  COR2X1 U1066 ( .A(n478), .B(n497), .Z(n1041) );
  COR2X1 U1067 ( .A(n518), .B(n535), .Z(n1042) );
  COR2X1 U1068 ( .A(n434), .B(n455), .Z(n1043) );
  CND2X1 U1069 ( .A(n498), .B(n517), .Z(n155) );
  COR2X1 U1070 ( .A(n600), .B(n613), .Z(n1045) );
  CND2X1 U1071 ( .A(n554), .B(n569), .Z(n178) );
  CND2X1 U1072 ( .A(n586), .B(n599), .Z(n188) );
  CND2X1 U1073 ( .A(n536), .B(n553), .Z(n172) );
  CND2X1 U1074 ( .A(n600), .B(n613), .Z(n200) );
  CND2X1 U1075 ( .A(n478), .B(n497), .Z(n152) );
  CND2X1 U1076 ( .A(n518), .B(n535), .Z(n167) );
  CND2X1 U1077 ( .A(n434), .B(n455), .Z(n132) );
  CND2X1 U1078 ( .A(n456), .B(n477), .Z(n141) );
  COND1XL U1079 ( .A(n236), .B(n232), .C(n233), .Z(n231) );
  COND1XL U1080 ( .A(n241), .B(n239), .C(n240), .Z(n238) );
  COND1XL U1081 ( .A(n1049), .B(n247), .C(n248), .Z(n246) );
  CANR1XL U1082 ( .A(n1050), .B(n246), .C(n243), .Z(n241) );
  CNR2X1 U1083 ( .A(n638), .B(n647), .Z(n213) );
  CNR2X1 U1084 ( .A(n666), .B(n673), .Z(n232) );
  CNR2X1 U1085 ( .A(n626), .B(n637), .Z(n210) );
  CENX1 U1086 ( .A(n80), .B(n234), .Z(product[10]) );
  COND1XL U1087 ( .A(n235), .B(n237), .C(n236), .Z(n234) );
  COR2X1 U1088 ( .A(n614), .B(n625), .Z(n1046) );
  COR2X1 U1089 ( .A(n648), .B(n657), .Z(n1048) );
  CND2X1 U1090 ( .A(n638), .B(n647), .Z(n214) );
  CND2X1 U1091 ( .A(n658), .B(n665), .Z(n227) );
  CND2X1 U1092 ( .A(n614), .B(n625), .Z(n205) );
  CND2X1 U1093 ( .A(n648), .B(n657), .Z(n222) );
  CENX1 U1094 ( .A(n83), .B(n246), .Z(product[7]) );
  CEOXL U1095 ( .A(n241), .B(n82), .Z(product[8]) );
  CND2X1 U1096 ( .A(n285), .B(n240), .Z(n82) );
  CEOX1 U1097 ( .A(n237), .B(n81), .Z(product[9]) );
  CNR2X1 U1098 ( .A(n690), .B(n693), .Z(n247) );
  CNR2X1 U1099 ( .A(n674), .B(n679), .Z(n235) );
  COAN1X1 U1100 ( .A(n251), .B(n253), .C(n252), .Z(n1049) );
  CNR2X1 U1101 ( .A(n680), .B(n685), .Z(n239) );
  COR2X1 U1102 ( .A(n686), .B(n689), .Z(n1050) );
  CND2X1 U1103 ( .A(n1051), .B(n89), .Z(n59) );
  CND2X1 U1104 ( .A(n305), .B(n291), .Z(n89) );
  CND2X1 U1105 ( .A(n674), .B(n679), .Z(n236) );
  CND2X1 U1106 ( .A(n686), .B(n689), .Z(n245) );
  COR2X1 U1107 ( .A(n305), .B(n291), .Z(n1051) );
  CENX1 U1108 ( .A(n86), .B(n258), .Z(product[4]) );
  CNR2X1 U1109 ( .A(n1062), .B(n16), .Z(n811) );
  CNR2X1 U1110 ( .A(n1063), .B(n15), .Z(n825) );
  CNR2X1 U1111 ( .A(n1057), .B(n24), .Z(n723) );
  CNR2X1 U1112 ( .A(n1062), .B(n18), .Z(n782) );
  CNR2X1 U1113 ( .A(n1063), .B(n17), .Z(n795) );
  CNR2X1 U1114 ( .A(n261), .B(n1052), .Z(n258) );
  CNR2X1 U1115 ( .A(n1055), .B(n1060), .Z(n933) );
  CNR2X1 U1116 ( .A(n1063), .B(n20), .Z(n756) );
  CNR2X1 U1117 ( .A(n694), .B(n695), .Z(n251) );
  CNR2X1 U1118 ( .A(n1057), .B(n23), .Z(n731) );
  CNR2X1 U1119 ( .A(n1057), .B(n20), .Z(n761) );
  CNR2X1 U1120 ( .A(n1065), .B(n962), .Z(n850) );
  CNR2X1 U1121 ( .A(n962), .B(n15), .Z(n818) );
  CNR2X1 U1122 ( .A(n1063), .B(n22), .Z(n735) );
  CNR2X1 U1123 ( .A(n1056), .B(n29), .Z(n699) );
  CNR2X1 U1124 ( .A(n1061), .B(n15), .Z(n827) );
  CNR2X1 U1125 ( .A(n1062), .B(n20), .Z(n757) );
  CNR2X1 U1126 ( .A(n1063), .B(n19), .Z(n768) );
  CNR2X1 U1127 ( .A(n1066), .B(n16), .Z(n807) );
  CNR2XL U1128 ( .A(n1064), .B(n19), .Z(n767) );
  CNR2X1 U1129 ( .A(n1062), .B(n1069), .Z(n876) );
  CNR2X1 U1130 ( .A(n1067), .B(n962), .Z(n849) );
  CNR2X1 U1131 ( .A(n1062), .B(n17), .Z(n796) );
  CNR2X1 U1132 ( .A(n1062), .B(n22), .Z(n736) );
  CNR2X1 U1133 ( .A(n1059), .B(n25), .Z(n715) );
  CNR2XL U1134 ( .A(n1064), .B(n23), .Z(n725) );
  CNR2X1 U1135 ( .A(n1062), .B(n21), .Z(n746) );
  CNR2X1 U1136 ( .A(n1057), .B(n25), .Z(n716) );
  CNR2X1 U1137 ( .A(n1062), .B(n24), .Z(n719) );
  CNR2X1 U1138 ( .A(n962), .B(n16), .Z(n803) );
  CNR2X1 U1139 ( .A(n1057), .B(n28), .Z(n701) );
  CNR2X1 U1140 ( .A(n1057), .B(n1064), .Z(n914) );
  CNR2X1 U1141 ( .A(n1059), .B(n1063), .Z(n919) );
  CNR2X1 U1142 ( .A(n1057), .B(n19), .Z(n773) );
  CNR2X1 U1143 ( .A(n1059), .B(n26), .Z(n709) );
  CNR2XL U1144 ( .A(n1064), .B(n21), .Z(n744) );
  CNR2X1 U1145 ( .A(n1063), .B(n16), .Z(n810) );
  CNR2X1 U1146 ( .A(n1054), .B(n22), .Z(n741) );
  CNR2X1 U1147 ( .A(n1063), .B(n21), .Z(n745) );
  CNR2X1 U1148 ( .A(n962), .B(n961), .Z(n832) );
  CNR2X1 U1149 ( .A(n1062), .B(n15), .Z(n826) );
  CNR2X1 U1150 ( .A(n1055), .B(n23), .Z(n732) );
  CNR2XL U1151 ( .A(n1064), .B(n16), .Z(n809) );
  CNR2X1 U1152 ( .A(n1063), .B(n18), .Z(n781) );
  CNR2XL U1153 ( .A(n1064), .B(n17), .Z(n794) );
  CNR2X1 U1154 ( .A(n1065), .B(n15), .Z(n823) );
  CNR2X1 U1155 ( .A(n1057), .B(n22), .Z(n740) );
  CNR2X1 U1156 ( .A(n1056), .B(n28), .Z(n702) );
  CNR2X1 U1157 ( .A(n1060), .B(n26), .Z(n708) );
  CNR2X1 U1158 ( .A(n961), .B(n15), .Z(n817) );
  CNR2X1 U1159 ( .A(n1057), .B(n21), .Z(n750) );
  CNR2X1 U1160 ( .A(n1065), .B(n961), .Z(n837) );
  CNR2X1 U1161 ( .A(n1060), .B(n19), .Z(n771) );
  CNR2X1 U1162 ( .A(n1069), .B(n1068), .Z(n871) );
  CNR2X1 U1163 ( .A(n1060), .B(n18), .Z(n784) );
  CNR2X1 U1164 ( .A(n1060), .B(n1068), .Z(n888) );
  CNR2X1 U1165 ( .A(n1062), .B(n962), .Z(n853) );
  CNR2X1 U1166 ( .A(n1061), .B(n961), .Z(n841) );
  CNR2X1 U1167 ( .A(n1061), .B(n1062), .Z(n922) );
  CNR2X1 U1168 ( .A(n1057), .B(n18), .Z(n786) );
  CNR2X1 U1169 ( .A(n1062), .B(n19), .Z(n769) );
  CNR2X1 U1170 ( .A(n1061), .B(n23), .Z(n728) );
  CNR2X1 U1171 ( .A(n1057), .B(n26), .Z(n710) );
  CNR2X1 U1172 ( .A(n1054), .B(n1067), .Z(n900) );
  CNR2X1 U1173 ( .A(n1063), .B(n961), .Z(n839) );
  CNR2X1 U1174 ( .A(n1060), .B(n17), .Z(n798) );
  CNR2X1 U1175 ( .A(n1056), .B(n26), .Z(n711) );
  CNR2X1 U1176 ( .A(n1061), .B(n1064), .Z(n911) );
  CNR2X1 U1177 ( .A(n1057), .B(n1068), .Z(n890) );
  CNR2X1 U1178 ( .A(n1063), .B(n963), .Z(n864) );
  CNR2X1 U1179 ( .A(n1056), .B(n27), .Z(n706) );
  CNR2X1 U1180 ( .A(n963), .B(n962), .Z(n846) );
  CNR2X1 U1181 ( .A(n1056), .B(n25), .Z(n717) );
  CNR2X1 U1182 ( .A(n1064), .B(n18), .Z(n780) );
  CNR2XL U1183 ( .A(n1064), .B(n22), .Z(n734) );
  CNR2X1 U1184 ( .A(n1057), .B(n1069), .Z(n880) );
  CNR2X1 U1185 ( .A(n1057), .B(n17), .Z(n800) );
  CNR2X1 U1186 ( .A(n1063), .B(n24), .Z(n718) );
  CND2X1 U1187 ( .A(n696), .B(n933), .Z(n257) );
  CEOX1 U1188 ( .A(n802), .B(n712), .Z(n304) );
  CNR2X1 U1189 ( .A(n961), .B(n16), .Z(n802) );
  CND2X1 U1190 ( .A(n694), .B(n695), .Z(n252) );
  COR2X1 U1191 ( .A(n696), .B(n933), .Z(n1053) );
  CNR2X1 U1192 ( .A(n1058), .B(n28), .Z(n700) );
  CNR2X1 U1193 ( .A(n1057), .B(n29), .Z(n698) );
  CNR2X1 U1194 ( .A(n962), .B(n17), .Z(n788) );
  CNR2X1 U1195 ( .A(n1057), .B(n1058), .Z(n934) );
  CNR2X1 U1196 ( .A(n1067), .B(n961), .Z(n836) );
  CNR2X1 U1197 ( .A(n1067), .B(n963), .Z(n861) );
  CNR2X1 U1198 ( .A(n1068), .B(n17), .Z(n791) );
  CNR2X1 U1199 ( .A(n1060), .B(n1063), .Z(n918) );
  CIVX2 U1200 ( .A(b[22]), .Z(n22) );
  CNR2X1 U1201 ( .A(n1056), .B(n30), .Z(n697) );
  CHA1XL U1202 ( .A(a[3]), .B(n929), .CO(n691), .S(n692) );
  CHA1XL U1203 ( .A(a[2]), .B(n934), .CO(n695), .S(n696) );
  CNR2XL U1204 ( .A(n1058), .B(n21), .Z(n749) );
  CNR2XL U1205 ( .A(n1058), .B(n24), .Z(n722) );
  CNR2X1 U1206 ( .A(n1059), .B(n17), .Z(n799) );
  CNR2X1 U1207 ( .A(n1058), .B(n23), .Z(n730) );
  CNR2X1 U1208 ( .A(n1058), .B(n18), .Z(n785) );
  CNR2X1 U1209 ( .A(n1059), .B(n19), .Z(n772) );
  CNR2X1 U1210 ( .A(n1058), .B(n20), .Z(n760) );
  CNR2X1 U1211 ( .A(n1059), .B(n22), .Z(n739) );
  CNR2X1 U1212 ( .A(n100), .B(n105), .Z(n98) );
  CNR2XL U1213 ( .A(n1065), .B(n22), .Z(n733) );
  CNR2XL U1214 ( .A(n1065), .B(n21), .Z(n743) );
  CNR2XL U1215 ( .A(n1065), .B(n20), .Z(n754) );
  CHA1XL U1216 ( .A(a[8]), .B(n886), .CO(n611), .S(n612) );
  CNR2X1 U1217 ( .A(n1065), .B(n16), .Z(n808) );
  CNR2X1 U1218 ( .A(n1065), .B(n17), .Z(n793) );
  CNR2X1 U1219 ( .A(n1065), .B(n19), .Z(n766) );
  CHA1XL U1220 ( .A(a[13]), .B(n821), .CO(n431), .S(n432) );
  CHA1XL U1221 ( .A(a[12]), .B(n836), .CO(n475), .S(n476) );
  CNR2XL U1222 ( .A(n1060), .B(n1065), .Z(n905) );
  CNR2X1 U1223 ( .A(n1062), .B(n1065), .Z(n903) );
  CNR2X1 U1224 ( .A(n1061), .B(n1065), .Z(n904) );
  CNR2X1 U1225 ( .A(n1063), .B(n1065), .Z(n902) );
  CNR2XL U1226 ( .A(n1059), .B(n1065), .Z(n906) );
  CHA1XL U1227 ( .A(a[4]), .B(n924), .CO(n683), .S(n684) );
  CIVX1 U1228 ( .A(b[1]), .Z(n1057) );
  CNR2X1 U1229 ( .A(n586), .B(n599), .Z(n187) );
  CHA1XL U1230 ( .A(a[9]), .B(n884), .CO(n583), .S(n584) );
  CNR2X1 U1231 ( .A(n1060), .B(n1066), .Z(n897) );
  CNR2XL U1232 ( .A(n1062), .B(n1066), .Z(n895) );
  CNR2XL U1233 ( .A(n1063), .B(n1066), .Z(n894) );
  CNR2X1 U1234 ( .A(n1064), .B(n1066), .Z(n893) );
  CNR2X1 U1235 ( .A(n1059), .B(n1066), .Z(n898) );
  CNR2X1 U1236 ( .A(n1065), .B(n1066), .Z(n892) );
  CNR2X1 U1237 ( .A(n1061), .B(n1066), .Z(n896) );
  COAN1X1 U1238 ( .A(n188), .B(n184), .C(n185), .Z(n181) );
  CNR2XL U1239 ( .A(n1070), .B(n19), .Z(n763) );
  CNR2X1 U1240 ( .A(n1070), .B(n962), .Z(n847) );
  CNR2X1 U1241 ( .A(n1070), .B(n963), .Z(n859) );
  CNR2X1 U1242 ( .A(n1070), .B(n15), .Z(n820) );
  CNR2XL U1243 ( .A(n1067), .B(n1070), .Z(n872) );
  CNR2X1 U1244 ( .A(n1070), .B(n961), .Z(n834) );
  CNR2XL U1245 ( .A(n1065), .B(n1070), .Z(n873) );
  CHA1XL U1246 ( .A(a[11]), .B(n861), .CO(n515), .S(n516) );
  CIVX1 U1247 ( .A(b[11]), .Z(n1069) );
  CNR2XL U1248 ( .A(n1065), .B(n1068), .Z(n883) );
  CNR2XL U1249 ( .A(n1062), .B(n1068), .Z(n886) );
  CNR2XL U1250 ( .A(n1068), .B(n962), .Z(n848) );
  CHA1XL U1251 ( .A(a[10]), .B(n882), .CO(n551), .S(n552) );
  CNR2XL U1252 ( .A(n1068), .B(n15), .Z(n821) );
  CNR2X1 U1253 ( .A(n1068), .B(n963), .Z(n860) );
  CNR2X1 U1254 ( .A(n1068), .B(n961), .Z(n835) );
  CHA1XL U1255 ( .A(a[6]), .B(n905), .CO(n655), .S(n656) );
  CIVXL U1256 ( .A(n174), .Z(n173) );
  COND1XL U1257 ( .A(n180), .B(n193), .C(n181), .Z(n179) );
  CNR2XL U1258 ( .A(n1064), .B(n1070), .Z(n874) );
  CNR2X1 U1259 ( .A(n1064), .B(n963), .Z(n863) );
  CNR2XL U1260 ( .A(n1064), .B(n1068), .Z(n884) );
  CNR2X1 U1261 ( .A(n1064), .B(n961), .Z(n838) );
  CHA1XL U1262 ( .A(a[7]), .B(n896), .CO(n635), .S(n636) );
  CNR2X1 U1263 ( .A(n1064), .B(n15), .Z(n824) );
  CNR2X1 U1264 ( .A(n1064), .B(n962), .Z(n851) );
  CEOXL U1265 ( .A(n63), .B(n118), .Z(product[27]) );
  CIVXL U1266 ( .A(n144), .Z(n146) );
  COND1XL U1267 ( .A(n143), .B(n160), .C(n144), .Z(n142) );
  CIVXL U1268 ( .A(\b[0] ), .Z(n1054) );
  CIVXL U1269 ( .A(\b[0] ), .Z(n1055) );
  CIVXL U1270 ( .A(\b[0] ), .Z(n1056) );
  CIVXL U1271 ( .A(b[2]), .Z(n1058) );
  CIVXL U1272 ( .A(b[2]), .Z(n1059) );
  CIVX2 U1273 ( .A(n94), .Z(n92) );
  CIVX2 U1274 ( .A(b[30]), .Z(n30) );
  CIVX2 U1275 ( .A(b[29]), .Z(n29) );
  CIVX2 U1276 ( .A(n251), .Z(n288) );
  CIVX2 U1277 ( .A(n247), .Z(n287) );
  CIVX2 U1278 ( .A(n239), .Z(n285) );
  CIVX2 U1279 ( .A(n235), .Z(n284) );
  CIVX2 U1280 ( .A(n232), .Z(n283) );
  CIVX2 U1281 ( .A(n213), .Z(n280) );
  CIVX2 U1282 ( .A(b[28]), .Z(n28) );
  CIVX2 U1283 ( .A(n210), .Z(n279) );
  CIVX2 U1284 ( .A(n177), .Z(n274) );
  CIVX2 U1285 ( .A(b[27]), .Z(n27) );
  CIVX2 U1286 ( .A(n116), .Z(n266) );
  CIVX2 U1287 ( .A(n105), .Z(n265) );
  CIVX2 U1288 ( .A(n100), .Z(n264) );
  CIVX2 U1289 ( .A(n257), .Z(n255) );
  CIVX2 U1290 ( .A(n245), .Z(n243) );
  CIVX2 U1291 ( .A(n238), .Z(n237) );
  CIVX2 U1292 ( .A(b[23]), .Z(n23) );
  CIVX2 U1293 ( .A(n229), .Z(n228) );
  CIVX2 U1294 ( .A(n227), .Z(n225) );
  CIVX2 U1295 ( .A(n222), .Z(n220) );
  CIVX2 U1296 ( .A(n216), .Z(n215) );
  CIVX2 U1297 ( .A(n207), .Z(n206) );
  CIVX2 U1298 ( .A(n205), .Z(n203) );
  CIVX2 U1299 ( .A(n200), .Z(n198) );
  CIVX2 U1300 ( .A(n194), .Z(n193) );
  CIVX2 U1301 ( .A(n187), .Z(n276) );
  CIVX2 U1302 ( .A(n184), .Z(n275) );
  CIVX2 U1303 ( .A(n172), .Z(n170) );
  CIVX2 U1304 ( .A(n167), .Z(n165) );
  CIVX2 U1305 ( .A(n155), .Z(n157) );
  CIVX2 U1306 ( .A(n154), .Z(n271) );
  CIVX2 U1307 ( .A(n143), .Z(n145) );
  CIVX2 U1308 ( .A(n141), .Z(n139) );
  CIVX2 U1309 ( .A(n132), .Z(n130) );
  CIVX2 U1310 ( .A(n124), .Z(n123) );
  CIVX2 U1311 ( .A(n122), .Z(n120) );
  CIVX2 U1312 ( .A(n121), .Z(n267) );
  CIVX2 U1313 ( .A(n111), .Z(n113) );
endmodule


module calc_DW_mult_uns_20 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n32, n36, n40, n44, n48, n52, n59, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n114, n115, n116, n117, n119, n121,
         n122, n123, n124, n128, n130, n131, n132, n133, n134, n135, n139,
         n141, n142, n143, n144, n146, n149, n150, n151, n152, n154, n156,
         n157, n158, n159, n160, n161, n162, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n177, n179, n180, n181,
         n182, n184, n187, n188, n189, n190, n192, n194, n195, n196, n197,
         n198, n199, n200, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n232,
         n234, n235, n236, n237, n240, n241, n242, n244, n246, n247, n250,
         n251, n253, n258, n260, n261, n262, n264, n266, n267, n268, n269,
         n270, n271, n272, n273, n275, n276, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n924, n949, n951, \b[0] , n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050;
  assign product[0] = \b[0] ;
  assign \b[0]  = b[0];

  CEO3X2 U298 ( .A(n297), .B(n280), .C(n295), .Z(n279) );
  CEO3X2 U299 ( .A(n299), .B(n282), .C(n281), .Z(n280) );
  CEO3X2 U300 ( .A(n284), .B(n283), .C(n301), .Z(n281) );
  CEO3X2 U301 ( .A(n286), .B(n303), .C(n285), .Z(n282) );
  CEO3X2 U302 ( .A(n287), .B(n307), .C(n305), .Z(n283) );
  CEO3X2 U303 ( .A(n291), .B(n289), .C(n288), .Z(n284) );
  CEO3X2 U304 ( .A(n311), .B(n290), .C(n309), .Z(n285) );
  CEO3X2 U305 ( .A(n317), .B(n315), .C(n313), .Z(n286) );
  CEO3X2 U306 ( .A(n730), .B(n319), .C(n292), .Z(n287) );
  CEO3X2 U307 ( .A(n751), .B(n713), .C(n691), .Z(n288) );
  CEO3X2 U308 ( .A(n776), .B(n700), .C(n686), .Z(n289) );
  CEO3X2 U309 ( .A(n763), .B(n695), .C(n706), .Z(n290) );
  CEO3X2 U310 ( .A(n740), .B(n790), .C(n721), .Z(n291) );
  CFA1X1 U312 ( .A(n298), .B(n296), .CI(n323), .CO(n293), .S(n294) );
  CFA1X1 U313 ( .A(n327), .B(n325), .CI(n300), .CO(n295), .S(n296) );
  CFA1X1 U314 ( .A(n304), .B(n302), .CI(n329), .CO(n297), .S(n298) );
  CFA1X1 U315 ( .A(n308), .B(n306), .CI(n331), .CO(n299), .S(n300) );
  CFA1X1 U316 ( .A(n310), .B(n333), .CI(n335), .CO(n301), .S(n302) );
  CFA1X1 U317 ( .A(n316), .B(n312), .CI(n314), .CO(n303), .S(n304) );
  CFA1X1 U318 ( .A(n337), .B(n318), .CI(n339), .CO(n305), .S(n306) );
  CFA1X1 U319 ( .A(n320), .B(n341), .CI(n343), .CO(n307), .S(n308) );
  CFA1X1 U320 ( .A(n741), .B(n345), .CI(n696), .CO(n309), .S(n310) );
  CFA1X1 U321 ( .A(n764), .B(n689), .CI(n722), .CO(n311), .S(n312) );
  CFA1X1 U322 ( .A(n752), .B(n707), .CI(n791), .CO(n313), .S(n314) );
  CFA1X1 U323 ( .A(n701), .B(n777), .CI(n731), .CO(n315), .S(n316) );
  CHA1X1 U325 ( .A(n687), .B(n714), .CO(n319), .S(n320) );
  CFA1X1 U326 ( .A(n326), .B(n324), .CI(n349), .CO(n321), .S(n322) );
  CFA1X1 U327 ( .A(n330), .B(n351), .CI(n328), .CO(n323), .S(n324) );
  CFA1X1 U328 ( .A(n332), .B(n353), .CI(n355), .CO(n325), .S(n326) );
  CFA1X1 U329 ( .A(n336), .B(n334), .CI(n357), .CO(n327), .S(n328) );
  CFA1X1 U330 ( .A(n340), .B(n359), .CI(n338), .CO(n329), .S(n330) );
  CFA1X1 U331 ( .A(n344), .B(n361), .CI(n342), .CO(n331), .S(n332) );
  CFA1X1 U332 ( .A(n367), .B(n363), .CI(n365), .CO(n333), .S(n334) );
  CFA1X1 U333 ( .A(n371), .B(n369), .CI(n346), .CO(n335), .S(n336) );
  CFA1X1 U334 ( .A(n753), .B(n702), .CI(n732), .CO(n337), .S(n338) );
  CFA1X1 U335 ( .A(n778), .B(n693), .CI(n715), .CO(n339), .S(n340) );
  CFA1X1 U336 ( .A(n697), .B(n806), .CI(n792), .CO(n341), .S(n342) );
  CFA1X1 U337 ( .A(n723), .B(n690), .CI(n765), .CO(n343), .S(n344) );
  CHA1X1 U338 ( .A(n742), .B(n708), .CO(n345), .S(n346) );
  CFA1X1 U339 ( .A(n352), .B(n350), .CI(n375), .CO(n347), .S(n348) );
  CFA1X1 U340 ( .A(n379), .B(n377), .CI(n354), .CO(n349), .S(n350) );
  CFA1X1 U341 ( .A(n381), .B(n356), .CI(n358), .CO(n351), .S(n352) );
  CFA1X1 U342 ( .A(n385), .B(n360), .CI(n383), .CO(n353), .S(n354) );
  CFA1X1 U343 ( .A(n387), .B(n362), .CI(n364), .CO(n355), .S(n356) );
  CFA1X1 U344 ( .A(n370), .B(n366), .CI(n368), .CO(n357), .S(n358) );
  CFA1X1 U345 ( .A(n393), .B(n389), .CI(n391), .CO(n359), .S(n360) );
  CFA1X1 U346 ( .A(n743), .B(n372), .CI(n395), .CO(n361), .S(n362) );
  CFA1X1 U347 ( .A(n766), .B(n698), .CI(n709), .CO(n363), .S(n364) );
  CFA1X1 U348 ( .A(n754), .B(n724), .CI(n820), .CO(n365), .S(n366) );
  CFA1X1 U349 ( .A(n716), .B(n793), .CI(n779), .CO(n367), .S(n368) );
  CFA1X1 U350 ( .A(n703), .B(n807), .CI(n733), .CO(n369), .S(n370) );
  CHA1X1 U351 ( .A(a[14]), .B(n694), .CO(n371), .S(n372) );
  CFA1X1 U352 ( .A(n378), .B(n376), .CI(n399), .CO(n373), .S(n374) );
  CFA1X1 U353 ( .A(n403), .B(n401), .CI(n380), .CO(n375), .S(n376) );
  CFA1X1 U354 ( .A(n405), .B(n382), .CI(n384), .CO(n377), .S(n378) );
  CFA1X1 U355 ( .A(n388), .B(n386), .CI(n407), .CO(n379), .S(n380) );
  CFA1X1 U356 ( .A(n392), .B(n409), .CI(n390), .CO(n381), .S(n382) );
  CFA1X1 U357 ( .A(n413), .B(n394), .CI(n411), .CO(n383), .S(n384) );
  CFA1X1 U358 ( .A(n396), .B(n415), .CI(n417), .CO(n385), .S(n386) );
  CFA1X1 U359 ( .A(n755), .B(n419), .CI(n734), .CO(n387), .S(n388) );
  CFA1X1 U360 ( .A(n780), .B(n704), .CI(n717), .CO(n389), .S(n390) );
  CFA1X1 U361 ( .A(n725), .B(n808), .CI(n794), .CO(n391), .S(n392) );
  CFA1X1 U362 ( .A(n699), .B(n710), .CI(n767), .CO(n393), .S(n394) );
  CHA1X1 U363 ( .A(n744), .B(n821), .CO(n395), .S(n396) );
  CFA1X1 U364 ( .A(n402), .B(n400), .CI(n423), .CO(n397), .S(n398) );
  CFA1X1 U365 ( .A(n427), .B(n425), .CI(n404), .CO(n399), .S(n400) );
  CFA1X1 U366 ( .A(n429), .B(n406), .CI(n408), .CO(n401), .S(n402) );
  CFA1X1 U367 ( .A(n412), .B(n410), .CI(n431), .CO(n403), .S(n404) );
  CFA1X1 U368 ( .A(n416), .B(n433), .CI(n414), .CO(n405), .S(n406) );
  CFA1X1 U369 ( .A(n437), .B(n418), .CI(n435), .CO(n407), .S(n408) );
  CFA1X1 U370 ( .A(n441), .B(n439), .CI(n420), .CO(n409), .S(n410) );
  CFA1X1 U371 ( .A(n768), .B(n711), .CI(n726), .CO(n411), .S(n412) );
  CFA1X1 U372 ( .A(n756), .B(n745), .CI(n834), .CO(n413), .S(n414) );
  CFA1X1 U373 ( .A(n735), .B(n795), .CI(n809), .CO(n415), .S(n416) );
  CFA1X1 U374 ( .A(n718), .B(n822), .CI(n781), .CO(n417), .S(n418) );
  CFA1X1 U376 ( .A(n426), .B(n424), .CI(n445), .CO(n421), .S(n422) );
  CFA1X1 U377 ( .A(n449), .B(n447), .CI(n428), .CO(n423), .S(n424) );
  CFA1X1 U378 ( .A(n451), .B(n430), .CI(n432), .CO(n425), .S(n426) );
  CFA1X1 U379 ( .A(n436), .B(n453), .CI(n434), .CO(n427), .S(n428) );
  CFA1X1 U380 ( .A(n455), .B(n438), .CI(n440), .CO(n429), .S(n430) );
  CFA1X1 U381 ( .A(n461), .B(n457), .CI(n459), .CO(n431), .S(n432) );
  CFA1X1 U382 ( .A(n757), .B(n442), .CI(n463), .CO(n433), .S(n434) );
  CFA1X1 U383 ( .A(n782), .B(n719), .CI(n736), .CO(n435), .S(n436) );
  CFA1X1 U384 ( .A(n727), .B(n835), .CI(n810), .CO(n437), .S(n438) );
  CFA1X1 U385 ( .A(n769), .B(n823), .CI(n796), .CO(n439), .S(n440) );
  CHA1X1 U386 ( .A(n746), .B(n712), .CO(n441), .S(n442) );
  CFA1X1 U387 ( .A(n448), .B(n446), .CI(n467), .CO(n443), .S(n444) );
  CFA1X1 U388 ( .A(n452), .B(n469), .CI(n450), .CO(n445), .S(n446) );
  CFA1X1 U389 ( .A(n473), .B(n471), .CI(n454), .CO(n447), .S(n448) );
  CFA1X1 U390 ( .A(n458), .B(n475), .CI(n456), .CO(n449), .S(n450) );
  CFA1X1 U391 ( .A(n477), .B(n460), .CI(n462), .CO(n451), .S(n452) );
  CFA1X1 U392 ( .A(n464), .B(n479), .CI(n481), .CO(n453), .S(n454) );
  CFA1X1 U393 ( .A(n797), .B(n483), .CI(n728), .CO(n455), .S(n456) );
  CFA1X1 U394 ( .A(n783), .B(n747), .CI(n847), .CO(n457), .S(n458) );
  CFA1X1 U395 ( .A(n758), .B(n770), .CI(n836), .CO(n459), .S(n460) );
  CFA1X1 U396 ( .A(n737), .B(n824), .CI(n811), .CO(n461), .S(n462) );
  CHA1X1 U397 ( .A(a[12]), .B(n720), .CO(n463), .S(n464) );
  CFA1X1 U398 ( .A(n470), .B(n468), .CI(n487), .CO(n465), .S(n466) );
  CFA1X1 U399 ( .A(n474), .B(n489), .CI(n472), .CO(n467), .S(n468) );
  CFA1X1 U400 ( .A(n493), .B(n491), .CI(n476), .CO(n469), .S(n470) );
  CFA1X1 U401 ( .A(n480), .B(n495), .CI(n478), .CO(n471), .S(n472) );
  CFA1X1 U402 ( .A(n501), .B(n482), .CI(n497), .CO(n473), .S(n474) );
  CFA1X1 U403 ( .A(n503), .B(n499), .CI(n484), .CO(n475), .S(n476) );
  CFA1X1 U404 ( .A(n784), .B(n738), .CI(n759), .CO(n477), .S(n478) );
  CFA1X1 U405 ( .A(n798), .B(n812), .CI(n837), .CO(n479), .S(n480) );
  CFA1X1 U406 ( .A(n771), .B(n729), .CI(n848), .CO(n481), .S(n482) );
  CHA1X1 U407 ( .A(n748), .B(n825), .CO(n483), .S(n484) );
  CFA1X1 U408 ( .A(n490), .B(n488), .CI(n507), .CO(n485), .S(n486) );
  CFA1X1 U409 ( .A(n494), .B(n509), .CI(n492), .CO(n487), .S(n488) );
  CFA1X1 U410 ( .A(n496), .B(n511), .CI(n513), .CO(n489), .S(n490) );
  CFA1X1 U411 ( .A(n502), .B(n498), .CI(n500), .CO(n491), .S(n492) );
  CFA1X1 U412 ( .A(n519), .B(n515), .CI(n517), .CO(n493), .S(n494) );
  CFA1X1 U413 ( .A(n772), .B(n504), .CI(n521), .CO(n495), .S(n496) );
  CFA1X1 U414 ( .A(n859), .B(n749), .CI(n849), .CO(n497), .S(n498) );
  CFA1X1 U416 ( .A(n760), .B(n799), .CI(n838), .CO(n501), .S(n502) );
  CHA1X1 U417 ( .A(n739), .B(n813), .CO(n503), .S(n504) );
  CFA1X1 U418 ( .A(n510), .B(n508), .CI(n525), .CO(n505), .S(n506) );
  CFA1X1 U419 ( .A(n529), .B(n527), .CI(n512), .CO(n507), .S(n508) );
  CFA1X1 U420 ( .A(n531), .B(n514), .CI(n516), .CO(n509), .S(n510) );
  CFA1X1 U421 ( .A(n533), .B(n518), .CI(n520), .CO(n511), .S(n512) );
  CFA1X1 U422 ( .A(n522), .B(n535), .CI(n537), .CO(n513), .S(n514) );
  CFA1X1 U423 ( .A(n860), .B(n539), .CI(n814), .CO(n515), .S(n516) );
  CFA1X1 U424 ( .A(n839), .B(n761), .CI(n786), .CO(n517), .S(n518) );
  CFA1X1 U425 ( .A(n800), .B(n850), .CI(n773), .CO(n519), .S(n520) );
  CHA1X1 U426 ( .A(n750), .B(n827), .CO(n521), .S(n522) );
  CFA1X1 U427 ( .A(n528), .B(n526), .CI(n543), .CO(n523), .S(n524) );
  CFA1X1 U428 ( .A(n532), .B(n545), .CI(n530), .CO(n525), .S(n526) );
  CFA1X1 U429 ( .A(n534), .B(n547), .CI(n549), .CO(n527), .S(n528) );
  CFA1X1 U430 ( .A(n551), .B(n536), .CI(n538), .CO(n529), .S(n530) );
  CFA1X1 U431 ( .A(n555), .B(n553), .CI(n540), .CO(n531), .S(n532) );
  CFA1X1 U432 ( .A(n840), .B(n828), .CI(n851), .CO(n533), .S(n534) );
  CFA1X1 U433 ( .A(n815), .B(n774), .CI(n870), .CO(n535), .S(n536) );
  CFA1X1 U434 ( .A(n787), .B(n801), .CI(n861), .CO(n537), .S(n538) );
  CHA1X1 U435 ( .A(a[10]), .B(n762), .CO(n539), .S(n540) );
  CFA1X1 U436 ( .A(n546), .B(n544), .CI(n559), .CO(n541), .S(n542) );
  CFA1X1 U437 ( .A(n563), .B(n548), .CI(n561), .CO(n543), .S(n544) );
  CFA1X1 U438 ( .A(n554), .B(n550), .CI(n552), .CO(n545), .S(n546) );
  CFA1X1 U439 ( .A(n569), .B(n565), .CI(n567), .CO(n547), .S(n548) );
  CFA1X1 U440 ( .A(n841), .B(n556), .CI(n571), .CO(n549), .S(n550) );
  CFA1X1 U441 ( .A(n862), .B(n788), .CI(n816), .CO(n551), .S(n552) );
  CFA1X1 U442 ( .A(n871), .B(n829), .CI(n802), .CO(n553), .S(n554) );
  CHA1X1 U443 ( .A(n775), .B(n852), .CO(n555), .S(n556) );
  CFA1X1 U444 ( .A(n562), .B(n560), .CI(n575), .CO(n557), .S(n558) );
  CFA1X1 U445 ( .A(n579), .B(n564), .CI(n577), .CO(n559), .S(n560) );
  CFA1X1 U446 ( .A(n570), .B(n566), .CI(n568), .CO(n561), .S(n562) );
  CFA1X1 U447 ( .A(n572), .B(n581), .CI(n583), .CO(n563), .S(n564) );
  CFA1X1 U448 ( .A(n872), .B(n585), .CI(n853), .CO(n565), .S(n566) );
  CFA1X1 U449 ( .A(n817), .B(n803), .CI(n880), .CO(n567), .S(n568) );
  CHA1X1 U451 ( .A(n789), .B(n863), .CO(n571), .S(n572) );
  CFA1X1 U452 ( .A(n578), .B(n576), .CI(n589), .CO(n573), .S(n574) );
  CFA1X1 U453 ( .A(n593), .B(n591), .CI(n580), .CO(n575), .S(n576) );
  CFA1X1 U454 ( .A(n597), .B(n582), .CI(n584), .CO(n577), .S(n578) );
  CFA1X1 U455 ( .A(n599), .B(n595), .CI(n586), .CO(n579), .S(n580) );
  CFA1X1 U456 ( .A(n881), .B(n818), .CI(n843), .CO(n581), .S(n582) );
  CFA1X1 U457 ( .A(n873), .B(n864), .CI(n854), .CO(n583), .S(n584) );
  CHA1X1 U458 ( .A(n804), .B(n831), .CO(n585), .S(n586) );
  CFA1X1 U459 ( .A(n592), .B(n590), .CI(n603), .CO(n587), .S(n588) );
  CFA1X1 U460 ( .A(n596), .B(n605), .CI(n594), .CO(n589), .S(n590) );
  CFA1X1 U461 ( .A(n609), .B(n598), .CI(n607), .CO(n591), .S(n592) );
  CFA1X1 U462 ( .A(n882), .B(n600), .CI(n611), .CO(n593), .S(n594) );
  CFA1X1 U463 ( .A(n865), .B(n855), .CI(n889), .CO(n595), .S(n596) );
  CFA1X1 U464 ( .A(n844), .B(n832), .CI(n874), .CO(n597), .S(n598) );
  CFA1X1 U466 ( .A(n606), .B(n604), .CI(n615), .CO(n601), .S(n602) );
  CFA1X1 U467 ( .A(n610), .B(n617), .CI(n608), .CO(n603), .S(n604) );
  CFA1X1 U468 ( .A(n612), .B(n621), .CI(n619), .CO(n605), .S(n606) );
  CFA1X1 U469 ( .A(n866), .B(n623), .CI(n845), .CO(n607), .S(n608) );
  CFA1X1 U470 ( .A(n856), .B(n883), .CI(n890), .CO(n609), .S(n610) );
  CHA1X1 U471 ( .A(n875), .B(n833), .CO(n611), .S(n612) );
  CFA1X1 U472 ( .A(n627), .B(n616), .CI(n618), .CO(n613), .S(n614) );
  CFA1X1 U473 ( .A(n622), .B(n629), .CI(n620), .CO(n615), .S(n616) );
  CFA1X1 U474 ( .A(n633), .B(n631), .CI(n624), .CO(n617), .S(n618) );
  CFA1X1 U475 ( .A(n867), .B(n876), .CI(n897), .CO(n619), .S(n620) );
  CFA1X1 U476 ( .A(n846), .B(n857), .CI(n891), .CO(n621), .S(n622) );
  CFA1X1 U478 ( .A(n630), .B(n628), .CI(n637), .CO(n625), .S(n626) );
  CFA1X1 U479 ( .A(n641), .B(n632), .CI(n639), .CO(n627), .S(n628) );
  CFA1X1 U480 ( .A(n868), .B(n634), .CI(n643), .CO(n629), .S(n630) );
  CFA1X1 U481 ( .A(n858), .B(n898), .CI(n885), .CO(n631), .S(n632) );
  CHA1X1 U482 ( .A(n877), .B(n892), .CO(n633), .S(n634) );
  CFA1X1 U483 ( .A(n640), .B(n638), .CI(n647), .CO(n635), .S(n636) );
  CFA1X1 U484 ( .A(n644), .B(n642), .CI(n649), .CO(n637), .S(n638) );
  CFA1X1 U485 ( .A(n899), .B(n651), .CI(n904), .CO(n639), .S(n640) );
  CFA1X1 U486 ( .A(n886), .B(n878), .CI(n893), .CO(n641), .S(n642) );
  CFA1X1 U488 ( .A(n650), .B(n648), .CI(n655), .CO(n645), .S(n646) );
  CFA1X1 U489 ( .A(n652), .B(n657), .CI(n659), .CO(n647), .S(n648) );
  CFA1X1 U490 ( .A(n905), .B(n887), .CI(n900), .CO(n649), .S(n650) );
  CHA1X1 U491 ( .A(n879), .B(n894), .CO(n651), .S(n652) );
  CFA1X1 U492 ( .A(n663), .B(n656), .CI(n658), .CO(n653), .S(n654) );
  CFA1X1 U493 ( .A(n910), .B(n660), .CI(n665), .CO(n655), .S(n656) );
  CFA1X1 U494 ( .A(n888), .B(n895), .CI(n906), .CO(n657), .S(n658) );
  CFA1X1 U496 ( .A(n671), .B(n664), .CI(n669), .CO(n661), .S(n662) );
  CFA1X1 U497 ( .A(n911), .B(n666), .CI(n902), .CO(n663), .S(n664) );
  CHA1X1 U498 ( .A(n896), .B(n907), .CO(n665), .S(n666) );
  CFA1X1 U499 ( .A(n675), .B(n670), .CI(n672), .CO(n667), .S(n668) );
  CFA1X1 U500 ( .A(n912), .B(n908), .CI(n915), .CO(n669), .S(n670) );
  CHA1X1 U501 ( .A(a[4]), .B(n903), .CO(n671), .S(n672) );
  CFA1X1 U502 ( .A(n913), .B(n679), .CI(n676), .CO(n673), .S(n674) );
  CHA1X1 U503 ( .A(n916), .B(n909), .CO(n675), .S(n676) );
  CFA1X1 U504 ( .A(n919), .B(n681), .CI(n917), .CO(n677), .S(n678) );
  CHA1X1 U506 ( .A(n918), .B(n920), .CO(n681), .S(n682) );
  CHA1X1 U507 ( .A(a[2]), .B(n921), .CO(n683), .S(n684) );
  CNR2X1 U796 ( .A(n32), .B(n951), .Z(n858) );
  COND1X1 U797 ( .A(n206), .B(n189), .C(n190), .Z(n188) );
  CHA1XL U798 ( .A(a[8]), .B(n819), .CO(n599), .S(n600) );
  CEOXL U799 ( .A(n80), .B(n218), .Z(product[11]) );
  CANR1XL U800 ( .A(n227), .B(n219), .C(n220), .Z(n218) );
  CENX1 U801 ( .A(n110), .B(n63), .Z(product[28]) );
  CIVX1 U802 ( .A(b[11]), .Z(n1047) );
  CIVX2 U803 ( .A(b[15]), .Z(n1050) );
  COR2X1 U804 ( .A(n924), .B(a[1]), .Z(n1025) );
  CNR2XL U805 ( .A(n949), .B(n16), .Z(n790) );
  CIVXL U806 ( .A(b[13]), .Z(n1049) );
  CIVXL U807 ( .A(b[13]), .Z(n1048) );
  CIVX2 U808 ( .A(b[2]), .Z(n36) );
  CFA1XL U809 ( .A(n692), .B(n805), .CI(a[15]), .CO(n317), .S(n318) );
  CIVX1 U810 ( .A(b[25]), .Z(n25) );
  CNR2XL U811 ( .A(n52), .B(n20), .Z(n740) );
  CNR2XL U812 ( .A(n19), .B(n52), .Z(n752) );
  CNR2XL U813 ( .A(n36), .B(n52), .Z(n877) );
  CNR2XL U814 ( .A(n17), .B(n52), .Z(n779) );
  CNR2XL U815 ( .A(n52), .B(n18), .Z(n765) );
  CNR2XL U816 ( .A(n1039), .B(n52), .Z(n878) );
  CNR2XL U817 ( .A(n1041), .B(n52), .Z(n876) );
  CNR2XL U818 ( .A(n48), .B(n52), .Z(n871) );
  CNR2XL U819 ( .A(n1042), .B(n52), .Z(n874) );
  CNR2XL U820 ( .A(n1047), .B(n52), .Z(n859) );
  CNR2XL U821 ( .A(n52), .B(n16), .Z(n794) );
  CNR2XL U822 ( .A(n1050), .B(n52), .Z(n809) );
  CNR2XL U823 ( .A(n1043), .B(n52), .Z(n872) );
  CIVXL U824 ( .A(b[23]), .Z(n23) );
  CIVXL U825 ( .A(b[17]), .Z(n17) );
  CENXL U826 ( .A(n1026), .B(n89), .Z(product[31]) );
  CNR2XL U827 ( .A(n1046), .B(n17), .Z(n780) );
  CIVXL U828 ( .A(b[16]), .Z(n16) );
  CNR2X1 U829 ( .A(n36), .B(n44), .Z(n907) );
  CANR1XL U830 ( .A(n207), .B(n215), .C(n208), .Z(n206) );
  CNR2XL U831 ( .A(n1050), .B(n36), .Z(n817) );
  CNR2XL U832 ( .A(n36), .B(n24), .Z(n710) );
  CND2X1 U833 ( .A(n1032), .B(n258), .Z(n132) );
  CNR2X1 U834 ( .A(n466), .B(n485), .Z(n143) );
  CNR2X1 U835 ( .A(n198), .B(n203), .Z(n196) );
  CANR1XL U836 ( .A(n1035), .B(n235), .C(n232), .Z(n230) );
  CANR1XL U837 ( .A(n247), .B(n1027), .C(n244), .Z(n242) );
  CNR2X1 U838 ( .A(n44), .B(n52), .Z(n873) );
  CNR2XL U839 ( .A(n1044), .B(n19), .Z(n755) );
  CNR2X1 U840 ( .A(n29), .B(n32), .Z(n687) );
  CNR2XL U841 ( .A(n40), .B(n52), .Z(n875) );
  CNR2X1 U842 ( .A(n1045), .B(n48), .Z(n880) );
  CNR2XL U843 ( .A(n1042), .B(n19), .Z(n757) );
  CNR2XL U844 ( .A(n1047), .B(n19), .Z(n751) );
  CNR2X1 U845 ( .A(n32), .B(n26), .Z(n699) );
  CIVX1 U846 ( .A(b[12]), .Z(n951) );
  CIVX1 U847 ( .A(b[14]), .Z(n949) );
  CIVX2 U848 ( .A(b[18]), .Z(n18) );
  CNR2X1 U849 ( .A(n1041), .B(n949), .Z(n830) );
  CNR2XL U850 ( .A(n1050), .B(n949), .Z(n805) );
  CND2XL U851 ( .A(n92), .B(n106), .Z(n90) );
  CND2XL U852 ( .A(n106), .B(n99), .Z(n97) );
  CND2IXL U853 ( .B(n111), .A(n112), .Z(n64) );
  CND2XL U854 ( .A(n99), .B(n102), .Z(n62) );
  CANR1X1 U855 ( .A(n146), .B(n1032), .C(n139), .Z(n133) );
  CIVX1 U856 ( .A(n141), .Z(n139) );
  COND1X1 U857 ( .A(n151), .B(n168), .C(n152), .Z(n150) );
  CND2XL U858 ( .A(n158), .B(n1031), .Z(n151) );
  CEOXL U859 ( .A(n70), .B(n162), .Z(product[21]) );
  CND2XL U860 ( .A(n260), .B(n161), .Z(n70) );
  CEOXL U861 ( .A(n69), .B(n157), .Z(product[22]) );
  CND2XL U862 ( .A(n1031), .B(n156), .Z(n69) );
  CEOXL U863 ( .A(n68), .B(n149), .Z(product[23]) );
  CND2XL U864 ( .A(n258), .B(n144), .Z(n68) );
  CND2XL U865 ( .A(n1030), .B(n194), .Z(n75) );
  CEOXL U866 ( .A(n74), .B(n187), .Z(product[17]) );
  CND2XL U867 ( .A(n264), .B(n182), .Z(n74) );
  CND2XL U868 ( .A(n1032), .B(n141), .Z(n67) );
  CND2XL U869 ( .A(n1029), .B(n130), .Z(n66) );
  CND2XL U870 ( .A(n1028), .B(n121), .Z(n65) );
  CND2XL U871 ( .A(n134), .B(n1029), .Z(n123) );
  CND2XL U872 ( .A(n261), .B(n166), .Z(n71) );
  CND2XL U873 ( .A(n348), .B(n373), .Z(n109) );
  CND2XL U874 ( .A(n294), .B(n321), .Z(n95) );
  CNR2XL U875 ( .A(n212), .B(n209), .Z(n207) );
  CANR1X1 U876 ( .A(n188), .B(n169), .C(n170), .Z(n168) );
  CNR2XL U877 ( .A(n174), .B(n171), .Z(n169) );
  COND1X1 U878 ( .A(n216), .B(n218), .C(n217), .Z(n215) );
  CND2XL U879 ( .A(n270), .B(n217), .Z(n80) );
  CND2XL U880 ( .A(n269), .B(n213), .Z(n79) );
  CND2XL U881 ( .A(n1033), .B(n179), .Z(n73) );
  CND2XL U882 ( .A(n262), .B(n172), .Z(n72) );
  CND2XL U883 ( .A(n267), .B(n204), .Z(n77) );
  CND2XL U884 ( .A(n1033), .B(n264), .Z(n174) );
  CIVXL U885 ( .A(n203), .Z(n267) );
  CIVXL U886 ( .A(n204), .Z(n202) );
  CNR2XL U887 ( .A(n221), .B(n224), .Z(n219) );
  CENX1 U888 ( .A(n279), .B(n293), .Z(n1026) );
  CND2XL U889 ( .A(n271), .B(n222), .Z(n81) );
  CND2XL U890 ( .A(n626), .B(n635), .Z(n210) );
  CND2XL U891 ( .A(n602), .B(n613), .Z(n199) );
  CND2XL U892 ( .A(n272), .B(n225), .Z(n82) );
  CND2XL U893 ( .A(n273), .B(n229), .Z(n83) );
  CEOXL U894 ( .A(n230), .B(n83), .Z(product[8]) );
  CND2XL U895 ( .A(n1035), .B(n234), .Z(n84) );
  CND2XL U896 ( .A(n276), .B(n241), .Z(n86) );
  CEOXL U897 ( .A(n242), .B(n86), .Z(product[5]) );
  CEOXL U898 ( .A(n1034), .B(n85), .Z(product[6]) );
  CND2XL U899 ( .A(n1027), .B(n246), .Z(n87) );
  CNR2XL U900 ( .A(n32), .B(n22), .Z(n729) );
  CNR2XL U901 ( .A(n1046), .B(n949), .Z(n824) );
  COR2X1 U902 ( .A(n684), .B(n922), .Z(n1027) );
  CNR2XL U903 ( .A(n44), .B(n24), .Z(n706) );
  CNR2XL U904 ( .A(n44), .B(n949), .Z(n827) );
  CNR2XL U905 ( .A(n32), .B(n20), .Z(n750) );
  CNR2XL U906 ( .A(n1041), .B(n1050), .Z(n816) );
  CNR2XL U907 ( .A(n1045), .B(n19), .Z(n753) );
  CNR2XL U908 ( .A(n1040), .B(n25), .Z(n702) );
  CNR2XL U909 ( .A(n1044), .B(n21), .Z(n732) );
  CNR2XL U910 ( .A(n1050), .B(n44), .Z(n813) );
  CNR2XL U911 ( .A(n21), .B(n32), .Z(n739) );
  CNR2XL U912 ( .A(n1046), .B(n1048), .Z(n837) );
  CNR2XL U913 ( .A(n1044), .B(n1050), .Z(n812) );
  CNR2XL U914 ( .A(n44), .B(n16), .Z(n798) );
  CNR2XL U915 ( .A(n1041), .B(n18), .Z(n772) );
  CNR2XL U916 ( .A(n1046), .B(n16), .Z(n795) );
  CNR2XL U917 ( .A(n1042), .B(n1045), .Z(n883) );
  CNR2XL U918 ( .A(n44), .B(n48), .Z(n890) );
  CNR2XL U919 ( .A(n21), .B(n44), .Z(n733) );
  CNR2XL U920 ( .A(n17), .B(n44), .Z(n783) );
  CNR2XL U921 ( .A(n1041), .B(n20), .Z(n747) );
  CNR2XL U922 ( .A(n1049), .B(n44), .Z(n840) );
  CNR2XL U923 ( .A(n1044), .B(n951), .Z(n851) );
  CNR2XL U924 ( .A(n44), .B(n22), .Z(n723) );
  CNR2XL U925 ( .A(n32), .B(n28), .Z(n690) );
  CNR2XL U926 ( .A(n1045), .B(n20), .Z(n741) );
  CNR2XL U927 ( .A(n1040), .B(n26), .Z(n696) );
  CNR2XL U928 ( .A(n1044), .B(n44), .Z(n897) );
  CNR2XL U929 ( .A(n1040), .B(n21), .Z(n736) );
  CNR2XL U930 ( .A(n1041), .B(n16), .Z(n801) );
  CNR2XL U931 ( .A(n1041), .B(n1044), .Z(n900) );
  CNR2XL U932 ( .A(n40), .B(n44), .Z(n905) );
  CNR2XL U933 ( .A(n1040), .B(n22), .Z(n726) );
  CNR2XL U934 ( .A(n1042), .B(n44), .Z(n904) );
  CNR2XL U935 ( .A(n1044), .B(n40), .Z(n899) );
  CNR2XL U936 ( .A(n1047), .B(n44), .Z(n863) );
  CNR2XL U937 ( .A(n17), .B(n32), .Z(n789) );
  CNR2XL U938 ( .A(n23), .B(n44), .Z(n714) );
  CNR2XL U939 ( .A(n32), .B(n949), .Z(n833) );
  CNR2XL U940 ( .A(n44), .B(n20), .Z(n744) );
  CNR2XL U941 ( .A(n1046), .B(n44), .Z(n882) );
  CNR2XL U942 ( .A(n1041), .B(n44), .Z(n906) );
  CNR2XL U943 ( .A(n1045), .B(n32), .Z(n888) );
  CNR2XL U944 ( .A(n44), .B(n18), .Z(n769) );
  CNR2XL U945 ( .A(n1041), .B(n19), .Z(n759) );
  CNR2XL U946 ( .A(n1045), .B(n18), .Z(n766) );
  CNR2XL U947 ( .A(n1040), .B(n24), .Z(n709) );
  CNR2XL U948 ( .A(n1041), .B(n1047), .Z(n866) );
  CNR2XL U949 ( .A(n19), .B(n44), .Z(n756) );
  CNR2XL U950 ( .A(n1039), .B(n32), .Z(n924) );
  CNR2XL U951 ( .A(n1040), .B(n951), .Z(n855) );
  CNR2XL U952 ( .A(n1046), .B(n52), .Z(n870) );
  CNR2XL U953 ( .A(n1040), .B(n23), .Z(n717) );
  CNR2XL U954 ( .A(n1049), .B(n32), .Z(n846) );
  CNR2XL U955 ( .A(n1046), .B(n1047), .Z(n860) );
  COR2XL U956 ( .A(n32), .B(n36), .Z(n1036) );
  CNR2XL U957 ( .A(n32), .B(n40), .Z(n918) );
  CNR2XL U958 ( .A(n32), .B(n52), .Z(n879) );
  CNR2XL U959 ( .A(n32), .B(n16), .Z(n804) );
  CNR2XL U960 ( .A(n1041), .B(n1042), .Z(n911) );
  CNR2XL U961 ( .A(n1042), .B(n1044), .Z(n898) );
  CNR2XL U962 ( .A(n1044), .B(n1048), .Z(n839) );
  CNR2XL U963 ( .A(n1041), .B(n48), .Z(n893) );
  CNR2XL U964 ( .A(n1046), .B(n36), .Z(n886) );
  CNR2XL U965 ( .A(n1040), .B(n1048), .Z(n843) );
  CNR2XL U966 ( .A(n1043), .B(n20), .Z(n743) );
  CNR2XL U967 ( .A(n1044), .B(n22), .Z(n722) );
  CNR2XL U968 ( .A(n32), .B(n48), .Z(n896) );
  CNR2XL U969 ( .A(n44), .B(n951), .Z(n852) );
  CNR2XL U970 ( .A(n32), .B(n18), .Z(n775) );
  CNR2XL U971 ( .A(n32), .B(n24), .Z(n712) );
  CNR2XL U972 ( .A(n1046), .B(n21), .Z(n730) );
  CND2XL U973 ( .A(n678), .B(n680), .Z(n237) );
  CNR2XL U974 ( .A(n1040), .B(n36), .Z(n919) );
  CNR2XL U975 ( .A(n1039), .B(n40), .Z(n917) );
  CNR2XL U976 ( .A(n1041), .B(n27), .Z(n691) );
  CEOXL U977 ( .A(n1036), .B(n250), .Z(product[3]) );
  CIVX1 U978 ( .A(b[4]), .Z(n40) );
  CIVX1 U979 ( .A(b[8]), .Z(n48) );
  CIVXL U980 ( .A(b[10]), .Z(n52) );
  CNR2XL U981 ( .A(n1049), .B(n40), .Z(n842) );
  CNR2XL U982 ( .A(n27), .B(n36), .Z(n692) );
  CNR2XL U983 ( .A(n1047), .B(n32), .Z(n869) );
  CNR2XL U984 ( .A(n1044), .B(n949), .Z(n826) );
  CNR2XL U985 ( .A(n17), .B(n40), .Z(n785) );
  CNR2XL U986 ( .A(n25), .B(n32), .Z(n705) );
  CIVXL U987 ( .A(b[19]), .Z(n19) );
  CNR2XL U988 ( .A(n1045), .B(n40), .Z(n884) );
  CIVXL U989 ( .A(b[20]), .Z(n20) );
  CIVXL U990 ( .A(b[22]), .Z(n22) );
  CNR2XL U991 ( .A(n23), .B(n32), .Z(n720) );
  CNR2XL U992 ( .A(n1042), .B(n32), .Z(n914) );
  CNR2XL U993 ( .A(n1044), .B(n32), .Z(n903) );
  CNR2XL U994 ( .A(n19), .B(n32), .Z(n762) );
  CNR2XL U995 ( .A(n1050), .B(n32), .Z(n819) );
  CNR2XL U996 ( .A(n27), .B(n32), .Z(n694) );
  CIVXL U997 ( .A(b[28]), .Z(n28) );
  CNR2XL U998 ( .A(n32), .B(n30), .Z(n685) );
  CAN2XL U999 ( .A(n1025), .B(n250), .Z(product[2]) );
  COND1XL U1000 ( .A(n112), .B(n108), .C(n109), .Z(n107) );
  CNR2X1 U1001 ( .A(n108), .B(n111), .Z(n106) );
  CANR1XL U1002 ( .A(n128), .B(n1028), .C(n119), .Z(n117) );
  CANR1XL U1003 ( .A(n99), .B(n107), .C(n100), .Z(n98) );
  CANR1XL U1004 ( .A(n107), .B(n92), .C(n93), .Z(n91) );
  COND1XL U1005 ( .A(n102), .B(n94), .C(n95), .Z(n93) );
  CND2X1 U1006 ( .A(n253), .B(n109), .Z(n63) );
  COND1XL U1007 ( .A(n111), .B(n59), .C(n112), .Z(n110) );
  CENX1 U1008 ( .A(n103), .B(n62), .Z(product[29]) );
  COND1XL U1009 ( .A(n104), .B(n59), .C(n105), .Z(n103) );
  CENX1 U1010 ( .A(n96), .B(n61), .Z(product[30]) );
  CND2X1 U1011 ( .A(n251), .B(n95), .Z(n61) );
  COND1XL U1012 ( .A(n97), .B(n59), .C(n98), .Z(n96) );
  CNR2X1 U1013 ( .A(n94), .B(n101), .Z(n92) );
  CANR1XL U1014 ( .A(n1031), .B(n159), .C(n154), .Z(n152) );
  CANR1X1 U1015 ( .A(n150), .B(n114), .C(n115), .Z(n59) );
  CNR2X1 U1016 ( .A(n116), .B(n132), .Z(n114) );
  COND1XL U1017 ( .A(n133), .B(n116), .C(n117), .Z(n115) );
  CND2X1 U1018 ( .A(n1028), .B(n1029), .Z(n116) );
  CND2X1 U1019 ( .A(n196), .B(n1030), .Z(n189) );
  CANR1XL U1020 ( .A(n1030), .B(n197), .C(n192), .Z(n190) );
  CNR2X1 U1021 ( .A(n374), .B(n397), .Z(n111) );
  COND1XL U1022 ( .A(n166), .B(n160), .C(n161), .Z(n159) );
  CNR2X1 U1023 ( .A(n348), .B(n373), .Z(n108) );
  CNR2X1 U1024 ( .A(n294), .B(n321), .Z(n94) );
  CANR1XL U1025 ( .A(n1029), .B(n135), .C(n128), .Z(n124) );
  CNR2X1 U1026 ( .A(n322), .B(n347), .Z(n101) );
  CENX1 U1027 ( .A(n142), .B(n67), .Z(product[24]) );
  COND1XL U1028 ( .A(n143), .B(n149), .C(n144), .Z(n142) );
  CENX1 U1029 ( .A(n131), .B(n66), .Z(product[25]) );
  COND1XL U1030 ( .A(n132), .B(n149), .C(n133), .Z(n131) );
  CENX1 U1031 ( .A(n122), .B(n65), .Z(product[26]) );
  COND1XL U1032 ( .A(n123), .B(n149), .C(n124), .Z(n122) );
  CENX1 U1033 ( .A(n167), .B(n71), .Z(product[20]) );
  CNR2X1 U1034 ( .A(n160), .B(n165), .Z(n158) );
  CEOX1 U1035 ( .A(n75), .B(n195), .Z(product[16]) );
  CANR1XL U1036 ( .A(n196), .B(n205), .C(n197), .Z(n195) );
  CANR1XL U1037 ( .A(n261), .B(n167), .C(n164), .Z(n162) );
  CANR1XL U1038 ( .A(n158), .B(n167), .C(n159), .Z(n157) );
  COR2X1 U1039 ( .A(n398), .B(n421), .Z(n1028) );
  CND2X1 U1040 ( .A(n322), .B(n347), .Z(n102) );
  CND2X1 U1041 ( .A(n374), .B(n397), .Z(n112) );
  CND2X1 U1042 ( .A(n398), .B(n421), .Z(n121) );
  COND1XL U1043 ( .A(n213), .B(n209), .C(n210), .Z(n208) );
  COND1XL U1044 ( .A(n171), .B(n175), .C(n172), .Z(n170) );
  CANR1XL U1045 ( .A(n184), .B(n1033), .C(n177), .Z(n175) );
  COND1XL U1046 ( .A(n204), .B(n198), .C(n199), .Z(n197) );
  CNR2X1 U1047 ( .A(n506), .B(n523), .Z(n160) );
  CNR2X1 U1048 ( .A(n524), .B(n541), .Z(n165) );
  COR2X1 U1049 ( .A(n422), .B(n443), .Z(n1029) );
  CENX1 U1050 ( .A(n211), .B(n78), .Z(product[13]) );
  CND2X1 U1051 ( .A(n268), .B(n210), .Z(n78) );
  COND1XL U1052 ( .A(n212), .B(n214), .C(n213), .Z(n211) );
  CENX1 U1053 ( .A(n205), .B(n77), .Z(product[14]) );
  CENX1 U1054 ( .A(n180), .B(n73), .Z(product[18]) );
  COND1XL U1055 ( .A(n181), .B(n187), .C(n182), .Z(n180) );
  CENX1 U1056 ( .A(n173), .B(n72), .Z(product[19]) );
  COND1XL U1057 ( .A(n174), .B(n187), .C(n175), .Z(n173) );
  CNR2X1 U1058 ( .A(n574), .B(n587), .Z(n181) );
  CEOX1 U1059 ( .A(n79), .B(n214), .Z(product[12]) );
  CEOX1 U1060 ( .A(n76), .B(n200), .Z(product[15]) );
  CND2X1 U1061 ( .A(n266), .B(n199), .Z(n76) );
  CANR1XL U1062 ( .A(n267), .B(n205), .C(n202), .Z(n200) );
  COR2X1 U1063 ( .A(n588), .B(n601), .Z(n1030) );
  COR2X1 U1064 ( .A(n486), .B(n505), .Z(n1031) );
  CND2X1 U1065 ( .A(n574), .B(n587), .Z(n182) );
  CND2X1 U1066 ( .A(n466), .B(n485), .Z(n144) );
  COR2X1 U1067 ( .A(n444), .B(n465), .Z(n1032) );
  CND2X1 U1068 ( .A(n524), .B(n541), .Z(n166) );
  CND2X1 U1069 ( .A(n422), .B(n443), .Z(n130) );
  CND2X1 U1070 ( .A(n588), .B(n601), .Z(n194) );
  CND2X1 U1071 ( .A(n486), .B(n505), .Z(n156) );
  CND2X1 U1072 ( .A(n444), .B(n465), .Z(n141) );
  CND2X1 U1073 ( .A(n506), .B(n523), .Z(n161) );
  COND1XL U1074 ( .A(n225), .B(n221), .C(n222), .Z(n220) );
  COND1XL U1075 ( .A(n230), .B(n228), .C(n229), .Z(n227) );
  CNR2X1 U1076 ( .A(n542), .B(n557), .Z(n171) );
  CNR2X1 U1077 ( .A(n626), .B(n635), .Z(n209) );
  CNR2X1 U1078 ( .A(n636), .B(n645), .Z(n212) );
  CNR2X1 U1079 ( .A(n602), .B(n613), .Z(n198) );
  CNR2X1 U1080 ( .A(n614), .B(n625), .Z(n203) );
  CENX1 U1081 ( .A(n81), .B(n223), .Z(product[10]) );
  COND1XL U1082 ( .A(n224), .B(n226), .C(n225), .Z(n223) );
  CNR2X1 U1083 ( .A(n646), .B(n653), .Z(n216) );
  COND1XL U1084 ( .A(n90), .B(n59), .C(n91), .Z(n89) );
  COR2X1 U1085 ( .A(n558), .B(n573), .Z(n1033) );
  CND2X1 U1086 ( .A(n614), .B(n625), .Z(n204) );
  CND2X1 U1087 ( .A(n636), .B(n645), .Z(n213) );
  CND2X1 U1088 ( .A(n558), .B(n573), .Z(n179) );
  CND2X1 U1089 ( .A(n646), .B(n653), .Z(n217) );
  CND2X1 U1090 ( .A(n542), .B(n557), .Z(n172) );
  CENX1 U1091 ( .A(n235), .B(n84), .Z(product[7]) );
  CEOX1 U1092 ( .A(n226), .B(n82), .Z(product[9]) );
  COND1XL U1093 ( .A(n1034), .B(n236), .C(n237), .Z(n235) );
  CNR2X1 U1094 ( .A(n662), .B(n667), .Z(n224) );
  CNR2X1 U1095 ( .A(n654), .B(n661), .Z(n221) );
  CNR2X1 U1096 ( .A(n668), .B(n673), .Z(n228) );
  COAN1X1 U1097 ( .A(n240), .B(n242), .C(n241), .Z(n1034) );
  CND2X1 U1098 ( .A(n662), .B(n667), .Z(n225) );
  CND2X1 U1099 ( .A(n674), .B(n677), .Z(n234) );
  CND2X1 U1100 ( .A(n654), .B(n661), .Z(n222) );
  CND2X1 U1101 ( .A(n668), .B(n673), .Z(n229) );
  COR2X1 U1102 ( .A(n674), .B(n677), .Z(n1035) );
  CND2X1 U1103 ( .A(n275), .B(n237), .Z(n85) );
  CNR2X1 U1104 ( .A(n949), .B(n52), .Z(n823) );
  CNR2X1 U1105 ( .A(n48), .B(n16), .Z(n796) );
  CNR2X1 U1106 ( .A(n1042), .B(n48), .Z(n891) );
  CNR2X1 U1107 ( .A(n1049), .B(n36), .Z(n844) );
  CNR2X1 U1108 ( .A(n23), .B(n40), .Z(n716) );
  CNR2X1 U1109 ( .A(n1047), .B(n16), .Z(n793) );
  CNR2X1 U1110 ( .A(n1042), .B(n17), .Z(n784) );
  CNR2X1 U1111 ( .A(n1043), .B(n16), .Z(n797) );
  CNR2X1 U1112 ( .A(n21), .B(n36), .Z(n737) );
  CNR2X1 U1113 ( .A(n1050), .B(n48), .Z(n811) );
  CNR2X1 U1114 ( .A(n1042), .B(n949), .Z(n828) );
  CNR2X1 U1115 ( .A(n1043), .B(n1047), .Z(n862) );
  CNR2X1 U1116 ( .A(n36), .B(n951), .Z(n856) );
  CNR2X1 U1117 ( .A(n1048), .B(n951), .Z(n834) );
  CNR2X1 U1118 ( .A(n1042), .B(n20), .Z(n745) );
  CNR2X1 U1119 ( .A(n1042), .B(n21), .Z(n734) );
  CNR2X1 U1120 ( .A(n682), .B(n683), .Z(n240) );
  CNR2X1 U1121 ( .A(n678), .B(n680), .Z(n236) );
  CNR2X1 U1122 ( .A(n25), .B(n36), .Z(n703) );
  CNR2X1 U1123 ( .A(n1050), .B(n951), .Z(n807) );
  CNR2X1 U1124 ( .A(n1048), .B(n48), .Z(n838) );
  CNR2X1 U1125 ( .A(n19), .B(n36), .Z(n760) );
  CNR2X1 U1126 ( .A(n1042), .B(n16), .Z(n799) );
  CNR2X1 U1127 ( .A(n17), .B(n951), .Z(n777) );
  CNR2X1 U1128 ( .A(n25), .B(n40), .Z(n701) );
  CNR2X1 U1129 ( .A(n21), .B(n48), .Z(n731) );
  CNR2X1 U1130 ( .A(n1043), .B(n17), .Z(n782) );
  CNR2X1 U1131 ( .A(n17), .B(n48), .Z(n781) );
  CNR2X1 U1132 ( .A(n23), .B(n36), .Z(n718) );
  CNR2X1 U1133 ( .A(n1047), .B(n949), .Z(n822) );
  CNR2X1 U1134 ( .A(n17), .B(n36), .Z(n787) );
  CNR2X1 U1135 ( .A(n1047), .B(n48), .Z(n861) );
  CNR2X1 U1136 ( .A(n1041), .B(n17), .Z(n786) );
  CNR2X1 U1137 ( .A(n1047), .B(n36), .Z(n867) );
  CNR2X1 U1138 ( .A(n1043), .B(n18), .Z(n768) );
  CNR2X1 U1139 ( .A(n1042), .B(n23), .Z(n715) );
  CNR2X1 U1140 ( .A(n1047), .B(n17), .Z(n778) );
  CNR2X1 U1141 ( .A(n951), .B(n52), .Z(n848) );
  CNR2X1 U1142 ( .A(n40), .B(n18), .Z(n771) );
  CNR2X1 U1143 ( .A(n1048), .B(n52), .Z(n836) );
  CNR2X1 U1144 ( .A(n19), .B(n40), .Z(n758) );
  CNR2X1 U1145 ( .A(n1042), .B(n18), .Z(n770) );
  CNR2X1 U1146 ( .A(n40), .B(n22), .Z(n725) );
  CNR2X1 U1147 ( .A(n1047), .B(n1050), .Z(n808) );
  CNR2X1 U1148 ( .A(n19), .B(n48), .Z(n754) );
  CNR2X1 U1149 ( .A(n1049), .B(n949), .Z(n820) );
  CNR2X1 U1150 ( .A(n1042), .B(n22), .Z(n724) );
  CNR2X1 U1151 ( .A(n40), .B(n951), .Z(n854) );
  CNR2X1 U1152 ( .A(n1042), .B(n1047), .Z(n864) );
  CNR2X1 U1153 ( .A(n951), .B(n16), .Z(n792) );
  CNR2X1 U1154 ( .A(n36), .B(n26), .Z(n697) );
  CNR2X1 U1155 ( .A(n1049), .B(n1050), .Z(n806) );
  CNR2X1 U1156 ( .A(n48), .B(n951), .Z(n850) );
  CNR2X1 U1157 ( .A(n40), .B(n16), .Z(n800) );
  CNR2X1 U1158 ( .A(n36), .B(n18), .Z(n773) );
  CNR2X1 U1159 ( .A(n1049), .B(n16), .Z(n791) );
  CNR2X1 U1160 ( .A(n1042), .B(n24), .Z(n707) );
  CNR2X1 U1161 ( .A(n951), .B(n949), .Z(n821) );
  CNR2X1 U1162 ( .A(n36), .B(n48), .Z(n894) );
  CNR2X1 U1163 ( .A(n36), .B(n949), .Z(n831) );
  CNR2X1 U1164 ( .A(n1040), .B(n1045), .Z(n885) );
  CNR2X1 U1165 ( .A(n21), .B(n40), .Z(n735) );
  CNR2X1 U1166 ( .A(n1050), .B(n40), .Z(n815) );
  CNR2X1 U1167 ( .A(n1042), .B(n951), .Z(n853) );
  CNR2X1 U1168 ( .A(n1047), .B(n40), .Z(n865) );
  CNR2X1 U1169 ( .A(n1043), .B(n48), .Z(n889) );
  CNR2X1 U1170 ( .A(n1047), .B(n951), .Z(n847) );
  CNR2X1 U1171 ( .A(n1042), .B(n1050), .Z(n814) );
  CNR2X1 U1172 ( .A(n40), .B(n949), .Z(n829) );
  CNR2X1 U1173 ( .A(n36), .B(n16), .Z(n802) );
  CNR2X1 U1174 ( .A(n36), .B(n40), .Z(n916) );
  CNR2X1 U1175 ( .A(n32), .B(n44), .Z(n909) );
  CNR2X1 U1176 ( .A(n48), .B(n20), .Z(n742) );
  CNR2X1 U1177 ( .A(n40), .B(n24), .Z(n708) );
  CNR2X1 U1178 ( .A(n48), .B(n949), .Z(n825) );
  CNR2X1 U1179 ( .A(n36), .B(n20), .Z(n748) );
  CNR2X1 U1180 ( .A(n1046), .B(n951), .Z(n849) );
  CNR2X1 U1181 ( .A(n1043), .B(n1045), .Z(n881) );
  CNR2X1 U1182 ( .A(n1042), .B(n40), .Z(n910) );
  CNR2X1 U1183 ( .A(n36), .B(n22), .Z(n727) );
  CNR2X1 U1184 ( .A(n1045), .B(n1050), .Z(n810) );
  CNR2X1 U1185 ( .A(n1047), .B(n1048), .Z(n835) );
  CNR2X1 U1186 ( .A(n1042), .B(n1048), .Z(n841) );
  CNR2X1 U1187 ( .A(n48), .B(n18), .Z(n767) );
  CNR2X1 U1188 ( .A(n1047), .B(n18), .Z(n764) );
  CNR2X1 U1189 ( .A(n1042), .B(n36), .Z(n912) );
  CNR2X1 U1190 ( .A(n1041), .B(n40), .Z(n915) );
  CNR2X1 U1191 ( .A(n40), .B(n48), .Z(n892) );
  CNR2X1 U1192 ( .A(n40), .B(n20), .Z(n746) );
  CEOX1 U1193 ( .A(n685), .B(n688), .Z(n292) );
  CNR2X1 U1194 ( .A(n1043), .B(n23), .Z(n713) );
  CNR2X1 U1195 ( .A(n40), .B(n26), .Z(n695) );
  CNR2X1 U1196 ( .A(n951), .B(n18), .Z(n763) );
  CNR2X1 U1197 ( .A(n48), .B(n22), .Z(n721) );
  CND2X1 U1198 ( .A(n682), .B(n683), .Z(n241) );
  CNR2X1 U1199 ( .A(n36), .B(n28), .Z(n688) );
  CNR2X1 U1200 ( .A(n1042), .B(n25), .Z(n700) );
  CNR2X1 U1201 ( .A(n1049), .B(n17), .Z(n776) );
  CIVX2 U1202 ( .A(\b[0] ), .Z(n32) );
  CNR2X1 U1203 ( .A(n1044), .B(n36), .Z(n901) );
  CNR2X1 U1204 ( .A(n1040), .B(n32), .Z(n921) );
  CIVX2 U1205 ( .A(b[6]), .Z(n44) );
  CHA1XL U1206 ( .A(a[6]), .B(n869), .CO(n643), .S(n644) );
  CEOXL U1207 ( .A(n64), .B(n59), .Z(product[27]) );
  CIVX1 U1208 ( .A(b[21]), .Z(n21) );
  CHA1XL U1209 ( .A(a[7]), .B(n884), .CO(n623), .S(n624) );
  CNR2X1 U1210 ( .A(n250), .B(n1036), .Z(n247) );
  CNR2X1 U1211 ( .A(n1038), .B(n48), .Z(n895) );
  CNR2XL U1212 ( .A(n1038), .B(n1044), .Z(n902) );
  CNR2X1 U1213 ( .A(n1038), .B(n44), .Z(n908) );
  CNR2X1 U1214 ( .A(n1039), .B(n1042), .Z(n913) );
  CNR2X1 U1215 ( .A(n1039), .B(n1040), .Z(n920) );
  CNR2X1 U1216 ( .A(n1039), .B(n36), .Z(n922) );
  CNR2X1 U1217 ( .A(n1038), .B(n16), .Z(n803) );
  CNR2X1 U1218 ( .A(n1038), .B(n17), .Z(n788) );
  CNR2X1 U1219 ( .A(n1038), .B(n18), .Z(n774) );
  CNR2X1 U1220 ( .A(n1038), .B(n19), .Z(n761) );
  CNR2X1 U1221 ( .A(n1038), .B(n20), .Z(n749) );
  CNR2X1 U1222 ( .A(n1038), .B(n21), .Z(n738) );
  CNR2X1 U1223 ( .A(n1038), .B(n22), .Z(n728) );
  CNR2X1 U1224 ( .A(n1038), .B(n23), .Z(n719) );
  CNR2X1 U1225 ( .A(n1038), .B(n24), .Z(n711) );
  CNR2X1 U1226 ( .A(n1039), .B(n25), .Z(n704) );
  CNR2X1 U1227 ( .A(n1039), .B(n26), .Z(n698) );
  CNR2X1 U1228 ( .A(n1039), .B(n27), .Z(n693) );
  CNR2X1 U1229 ( .A(n1039), .B(n28), .Z(n689) );
  CNR2X1 U1230 ( .A(n1039), .B(n29), .Z(n686) );
  CNR2XL U1231 ( .A(n1038), .B(n1050), .Z(n818) );
  CNR2X1 U1232 ( .A(n1038), .B(n949), .Z(n832) );
  CNR2X1 U1233 ( .A(n1038), .B(n1048), .Z(n845) );
  CNR2X1 U1234 ( .A(n1039), .B(n951), .Z(n857) );
  CNR2XL U1235 ( .A(n1039), .B(n1047), .Z(n868) );
  CNR2XL U1236 ( .A(n1039), .B(n1045), .Z(n887) );
  CENX1 U1237 ( .A(n87), .B(n247), .Z(product[4]) );
  CND2X1 U1238 ( .A(n684), .B(n922), .Z(n246) );
  CND2XL U1239 ( .A(n924), .B(a[1]), .Z(n250) );
  CIVX1 U1240 ( .A(b[5]), .Z(n1042) );
  CFA1XL U1241 ( .A(a[9]), .B(n830), .CI(n842), .CO(n569), .S(n570) );
  CHA1XL U1242 ( .A(a[3]), .B(n914), .CO(n679), .S(n680) );
  CFA1XL U1243 ( .A(a[11]), .B(n826), .CI(n785), .CO(n499), .S(n500) );
  CHA1XL U1244 ( .A(n705), .B(a[13]), .CO(n419), .S(n420) );
  CHA1XL U1245 ( .A(a[5]), .B(n901), .CO(n659), .S(n660) );
  CIVXL U1246 ( .A(b[1]), .Z(n1038) );
  CIVXL U1247 ( .A(b[1]), .Z(n1039) );
  CIVXL U1248 ( .A(b[3]), .Z(n1040) );
  CIVXL U1249 ( .A(b[3]), .Z(n1041) );
  CIVXL U1250 ( .A(b[7]), .Z(n1043) );
  CIVXL U1251 ( .A(b[7]), .Z(n1044) );
  CIVXL U1252 ( .A(b[9]), .Z(n1045) );
  CIVXL U1253 ( .A(b[9]), .Z(n1046) );
  CIVX2 U1254 ( .A(b[30]), .Z(n30) );
  CIVX2 U1255 ( .A(b[29]), .Z(n29) );
  CIVX2 U1256 ( .A(n240), .Z(n276) );
  CIVX2 U1257 ( .A(n236), .Z(n275) );
  CIVX2 U1258 ( .A(n228), .Z(n273) );
  CIVX2 U1259 ( .A(n224), .Z(n272) );
  CIVX2 U1260 ( .A(n221), .Z(n271) );
  CIVX2 U1261 ( .A(n216), .Z(n270) );
  CIVX2 U1262 ( .A(b[27]), .Z(n27) );
  CIVX2 U1263 ( .A(n212), .Z(n269) );
  CIVX2 U1264 ( .A(n209), .Z(n268) );
  CIVX2 U1265 ( .A(n198), .Z(n266) );
  CIVX2 U1266 ( .A(n171), .Z(n262) );
  CIVX2 U1267 ( .A(n160), .Z(n260) );
  CIVX2 U1268 ( .A(b[26]), .Z(n26) );
  CIVX2 U1269 ( .A(n108), .Z(n253) );
  CIVX2 U1270 ( .A(n101), .Z(n99) );
  CIVX2 U1271 ( .A(n94), .Z(n251) );
  CIVX2 U1272 ( .A(n246), .Z(n244) );
  CIVX2 U1273 ( .A(b[24]), .Z(n24) );
  CIVX2 U1274 ( .A(n234), .Z(n232) );
  CIVX2 U1275 ( .A(n227), .Z(n226) );
  CIVX2 U1276 ( .A(n215), .Z(n214) );
  CIVX2 U1277 ( .A(n206), .Z(n205) );
  CIVX2 U1278 ( .A(n194), .Z(n192) );
  CIVX2 U1279 ( .A(n188), .Z(n187) );
  CIVX2 U1280 ( .A(n182), .Z(n184) );
  CIVX2 U1281 ( .A(n181), .Z(n264) );
  CIVX2 U1282 ( .A(n179), .Z(n177) );
  CIVX2 U1283 ( .A(n168), .Z(n167) );
  CIVX2 U1284 ( .A(n166), .Z(n164) );
  CIVX2 U1285 ( .A(n165), .Z(n261) );
  CIVX2 U1286 ( .A(n156), .Z(n154) );
  CIVX2 U1287 ( .A(n150), .Z(n149) );
  CIVX2 U1288 ( .A(n144), .Z(n146) );
  CIVX2 U1289 ( .A(n143), .Z(n258) );
  CIVX2 U1290 ( .A(n133), .Z(n135) );
  CIVX2 U1291 ( .A(n132), .Z(n134) );
  CIVX2 U1292 ( .A(n130), .Z(n128) );
  CIVX2 U1293 ( .A(n121), .Z(n119) );
  CIVX2 U1294 ( .A(n107), .Z(n105) );
  CIVX2 U1295 ( .A(n106), .Z(n104) );
  CIVX2 U1296 ( .A(n102), .Z(n100) );
endmodule


module calc_DW_mult_uns_21 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n32, n36, n40, n44, n48, n52, n59, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n114, n115, n116, n117, n119, n121,
         n122, n123, n124, n128, n130, n131, n132, n133, n134, n135, n139,
         n141, n142, n143, n144, n146, n149, n150, n151, n152, n154, n156,
         n157, n158, n159, n160, n161, n162, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n177, n179, n180, n181,
         n182, n184, n187, n188, n189, n190, n192, n194, n195, n196, n197,
         n198, n199, n200, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n232,
         n234, n235, n236, n237, n240, n241, n242, n244, n246, n247, n250,
         n251, n253, n258, n260, n261, n262, n264, n266, n267, n268, n269,
         n270, n271, n272, n273, n275, n276, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n924, n949, n951, \b[0] , n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048;
  assign product[0] = \b[0] ;
  assign \b[0]  = b[0];

  CANR1X1 U164 ( .A(n188), .B(n169), .C(n170), .Z(n168) );
  CEO3X2 U298 ( .A(n297), .B(n280), .C(n295), .Z(n279) );
  CEO3X2 U299 ( .A(n299), .B(n282), .C(n281), .Z(n280) );
  CEO3X2 U300 ( .A(n284), .B(n283), .C(n301), .Z(n281) );
  CEO3X2 U301 ( .A(n286), .B(n303), .C(n285), .Z(n282) );
  CEO3X2 U302 ( .A(n287), .B(n307), .C(n305), .Z(n283) );
  CEO3X2 U303 ( .A(n291), .B(n289), .C(n288), .Z(n284) );
  CEO3X2 U304 ( .A(n311), .B(n290), .C(n309), .Z(n285) );
  CEO3X2 U305 ( .A(n317), .B(n315), .C(n313), .Z(n286) );
  CEO3X2 U306 ( .A(n730), .B(n319), .C(n292), .Z(n287) );
  CEO3X2 U307 ( .A(n751), .B(n713), .C(n691), .Z(n288) );
  CEO3X2 U308 ( .A(n776), .B(n700), .C(n686), .Z(n289) );
  CEO3X2 U309 ( .A(n763), .B(n695), .C(n706), .Z(n290) );
  CEO3X2 U310 ( .A(n740), .B(n790), .C(n721), .Z(n291) );
  CFA1X1 U312 ( .A(n298), .B(n296), .CI(n323), .CO(n293), .S(n294) );
  CFA1X1 U313 ( .A(n327), .B(n325), .CI(n300), .CO(n295), .S(n296) );
  CFA1X1 U314 ( .A(n304), .B(n302), .CI(n329), .CO(n297), .S(n298) );
  CFA1X1 U315 ( .A(n308), .B(n306), .CI(n331), .CO(n299), .S(n300) );
  CFA1X1 U316 ( .A(n310), .B(n333), .CI(n335), .CO(n301), .S(n302) );
  CFA1X1 U317 ( .A(n316), .B(n312), .CI(n314), .CO(n303), .S(n304) );
  CFA1X1 U318 ( .A(n337), .B(n318), .CI(n339), .CO(n305), .S(n306) );
  CFA1X1 U319 ( .A(n320), .B(n341), .CI(n343), .CO(n307), .S(n308) );
  CFA1X1 U320 ( .A(n741), .B(n345), .CI(n696), .CO(n309), .S(n310) );
  CFA1X1 U321 ( .A(n764), .B(n689), .CI(n722), .CO(n311), .S(n312) );
  CFA1X1 U322 ( .A(n752), .B(n707), .CI(n791), .CO(n313), .S(n314) );
  CFA1X1 U323 ( .A(n701), .B(n777), .CI(n731), .CO(n315), .S(n316) );
  CFA1X1 U324 ( .A(n692), .B(n805), .CI(a[15]), .CO(n317), .S(n318) );
  CHA1X1 U325 ( .A(n687), .B(n714), .CO(n319), .S(n320) );
  CFA1X1 U326 ( .A(n326), .B(n324), .CI(n349), .CO(n321), .S(n322) );
  CFA1X1 U327 ( .A(n330), .B(n351), .CI(n328), .CO(n323), .S(n324) );
  CFA1X1 U328 ( .A(n332), .B(n353), .CI(n355), .CO(n325), .S(n326) );
  CFA1X1 U329 ( .A(n336), .B(n334), .CI(n357), .CO(n327), .S(n328) );
  CFA1X1 U330 ( .A(n340), .B(n359), .CI(n338), .CO(n329), .S(n330) );
  CFA1X1 U331 ( .A(n344), .B(n361), .CI(n342), .CO(n331), .S(n332) );
  CFA1X1 U332 ( .A(n367), .B(n363), .CI(n365), .CO(n333), .S(n334) );
  CFA1X1 U333 ( .A(n371), .B(n369), .CI(n346), .CO(n335), .S(n336) );
  CFA1X1 U334 ( .A(n753), .B(n702), .CI(n732), .CO(n337), .S(n338) );
  CFA1X1 U335 ( .A(n778), .B(n693), .CI(n715), .CO(n339), .S(n340) );
  CFA1X1 U336 ( .A(n697), .B(n806), .CI(n792), .CO(n341), .S(n342) );
  CFA1X1 U337 ( .A(n723), .B(n690), .CI(n765), .CO(n343), .S(n344) );
  CHA1X1 U338 ( .A(n742), .B(n708), .CO(n345), .S(n346) );
  CFA1X1 U339 ( .A(n352), .B(n350), .CI(n375), .CO(n347), .S(n348) );
  CFA1X1 U340 ( .A(n379), .B(n377), .CI(n354), .CO(n349), .S(n350) );
  CFA1X1 U341 ( .A(n381), .B(n356), .CI(n358), .CO(n351), .S(n352) );
  CFA1X1 U342 ( .A(n385), .B(n360), .CI(n383), .CO(n353), .S(n354) );
  CFA1X1 U343 ( .A(n387), .B(n362), .CI(n364), .CO(n355), .S(n356) );
  CFA1X1 U344 ( .A(n370), .B(n366), .CI(n368), .CO(n357), .S(n358) );
  CFA1X1 U345 ( .A(n393), .B(n389), .CI(n391), .CO(n359), .S(n360) );
  CFA1X1 U346 ( .A(n743), .B(n372), .CI(n395), .CO(n361), .S(n362) );
  CFA1X1 U347 ( .A(n766), .B(n698), .CI(n709), .CO(n363), .S(n364) );
  CFA1X1 U348 ( .A(n754), .B(n724), .CI(n820), .CO(n365), .S(n366) );
  CFA1X1 U349 ( .A(n716), .B(n793), .CI(n779), .CO(n367), .S(n368) );
  CFA1X1 U350 ( .A(n703), .B(n807), .CI(n733), .CO(n369), .S(n370) );
  CHA1X1 U351 ( .A(a[14]), .B(n694), .CO(n371), .S(n372) );
  CFA1X1 U352 ( .A(n378), .B(n376), .CI(n399), .CO(n373), .S(n374) );
  CFA1X1 U353 ( .A(n403), .B(n401), .CI(n380), .CO(n375), .S(n376) );
  CFA1X1 U354 ( .A(n405), .B(n382), .CI(n384), .CO(n377), .S(n378) );
  CFA1X1 U355 ( .A(n388), .B(n386), .CI(n407), .CO(n379), .S(n380) );
  CFA1X1 U356 ( .A(n392), .B(n409), .CI(n390), .CO(n381), .S(n382) );
  CFA1X1 U357 ( .A(n413), .B(n394), .CI(n411), .CO(n383), .S(n384) );
  CFA1X1 U358 ( .A(n396), .B(n415), .CI(n417), .CO(n385), .S(n386) );
  CFA1X1 U359 ( .A(n755), .B(n419), .CI(n734), .CO(n387), .S(n388) );
  CFA1X1 U360 ( .A(n780), .B(n704), .CI(n717), .CO(n389), .S(n390) );
  CFA1X1 U361 ( .A(n725), .B(n808), .CI(n794), .CO(n391), .S(n392) );
  CFA1X1 U362 ( .A(n699), .B(n710), .CI(n767), .CO(n393), .S(n394) );
  CHA1X1 U363 ( .A(n744), .B(n821), .CO(n395), .S(n396) );
  CFA1X1 U364 ( .A(n402), .B(n400), .CI(n423), .CO(n397), .S(n398) );
  CFA1X1 U365 ( .A(n427), .B(n425), .CI(n404), .CO(n399), .S(n400) );
  CFA1X1 U366 ( .A(n429), .B(n406), .CI(n408), .CO(n401), .S(n402) );
  CFA1X1 U367 ( .A(n412), .B(n410), .CI(n431), .CO(n403), .S(n404) );
  CFA1X1 U368 ( .A(n416), .B(n433), .CI(n414), .CO(n405), .S(n406) );
  CFA1X1 U369 ( .A(n437), .B(n418), .CI(n435), .CO(n407), .S(n408) );
  CFA1X1 U370 ( .A(n441), .B(n439), .CI(n420), .CO(n409), .S(n410) );
  CFA1X1 U371 ( .A(n768), .B(n711), .CI(n726), .CO(n411), .S(n412) );
  CFA1X1 U372 ( .A(n756), .B(n745), .CI(n834), .CO(n413), .S(n414) );
  CFA1X1 U373 ( .A(n735), .B(n795), .CI(n809), .CO(n415), .S(n416) );
  CFA1X1 U374 ( .A(n718), .B(n822), .CI(n781), .CO(n417), .S(n418) );
  CFA1X1 U376 ( .A(n426), .B(n424), .CI(n445), .CO(n421), .S(n422) );
  CFA1X1 U377 ( .A(n449), .B(n447), .CI(n428), .CO(n423), .S(n424) );
  CFA1X1 U378 ( .A(n451), .B(n430), .CI(n432), .CO(n425), .S(n426) );
  CFA1X1 U379 ( .A(n436), .B(n453), .CI(n434), .CO(n427), .S(n428) );
  CFA1X1 U380 ( .A(n455), .B(n438), .CI(n440), .CO(n429), .S(n430) );
  CFA1X1 U381 ( .A(n461), .B(n457), .CI(n459), .CO(n431), .S(n432) );
  CFA1X1 U382 ( .A(n757), .B(n442), .CI(n463), .CO(n433), .S(n434) );
  CFA1X1 U383 ( .A(n782), .B(n719), .CI(n736), .CO(n435), .S(n436) );
  CFA1X1 U384 ( .A(n727), .B(n835), .CI(n810), .CO(n437), .S(n438) );
  CFA1X1 U385 ( .A(n769), .B(n823), .CI(n796), .CO(n439), .S(n440) );
  CHA1X1 U386 ( .A(n746), .B(n712), .CO(n441), .S(n442) );
  CFA1X1 U387 ( .A(n448), .B(n446), .CI(n467), .CO(n443), .S(n444) );
  CFA1X1 U388 ( .A(n452), .B(n469), .CI(n450), .CO(n445), .S(n446) );
  CFA1X1 U389 ( .A(n473), .B(n471), .CI(n454), .CO(n447), .S(n448) );
  CFA1X1 U390 ( .A(n458), .B(n475), .CI(n456), .CO(n449), .S(n450) );
  CFA1X1 U391 ( .A(n477), .B(n460), .CI(n462), .CO(n451), .S(n452) );
  CFA1X1 U392 ( .A(n464), .B(n479), .CI(n481), .CO(n453), .S(n454) );
  CFA1X1 U393 ( .A(n797), .B(n483), .CI(n728), .CO(n455), .S(n456) );
  CFA1X1 U394 ( .A(n783), .B(n747), .CI(n847), .CO(n457), .S(n458) );
  CFA1X1 U395 ( .A(n758), .B(n770), .CI(n836), .CO(n459), .S(n460) );
  CFA1X1 U396 ( .A(n737), .B(n824), .CI(n811), .CO(n461), .S(n462) );
  CHA1X1 U397 ( .A(a[12]), .B(n720), .CO(n463), .S(n464) );
  CFA1X1 U398 ( .A(n470), .B(n468), .CI(n487), .CO(n465), .S(n466) );
  CFA1X1 U399 ( .A(n474), .B(n489), .CI(n472), .CO(n467), .S(n468) );
  CFA1X1 U400 ( .A(n493), .B(n491), .CI(n476), .CO(n469), .S(n470) );
  CFA1X1 U401 ( .A(n480), .B(n495), .CI(n478), .CO(n471), .S(n472) );
  CFA1X1 U402 ( .A(n501), .B(n482), .CI(n497), .CO(n473), .S(n474) );
  CFA1X1 U403 ( .A(n503), .B(n499), .CI(n484), .CO(n475), .S(n476) );
  CFA1X1 U404 ( .A(n784), .B(n738), .CI(n759), .CO(n477), .S(n478) );
  CFA1X1 U405 ( .A(n798), .B(n812), .CI(n837), .CO(n479), .S(n480) );
  CFA1X1 U406 ( .A(n771), .B(n729), .CI(n848), .CO(n481), .S(n482) );
  CHA1X1 U407 ( .A(n748), .B(n825), .CO(n483), .S(n484) );
  CFA1X1 U408 ( .A(n490), .B(n488), .CI(n507), .CO(n485), .S(n486) );
  CFA1X1 U409 ( .A(n494), .B(n509), .CI(n492), .CO(n487), .S(n488) );
  CFA1X1 U410 ( .A(n496), .B(n511), .CI(n513), .CO(n489), .S(n490) );
  CFA1X1 U411 ( .A(n502), .B(n498), .CI(n500), .CO(n491), .S(n492) );
  CFA1X1 U412 ( .A(n519), .B(n515), .CI(n517), .CO(n493), .S(n494) );
  CFA1X1 U413 ( .A(n772), .B(n504), .CI(n521), .CO(n495), .S(n496) );
  CFA1X1 U414 ( .A(n859), .B(n749), .CI(n849), .CO(n497), .S(n498) );
  CFA1X1 U416 ( .A(n760), .B(n799), .CI(n838), .CO(n501), .S(n502) );
  CHA1X1 U417 ( .A(n739), .B(n813), .CO(n503), .S(n504) );
  CFA1X1 U418 ( .A(n510), .B(n508), .CI(n525), .CO(n505), .S(n506) );
  CFA1X1 U419 ( .A(n529), .B(n527), .CI(n512), .CO(n507), .S(n508) );
  CFA1X1 U420 ( .A(n531), .B(n514), .CI(n516), .CO(n509), .S(n510) );
  CFA1X1 U421 ( .A(n533), .B(n518), .CI(n520), .CO(n511), .S(n512) );
  CFA1X1 U422 ( .A(n522), .B(n535), .CI(n537), .CO(n513), .S(n514) );
  CFA1X1 U423 ( .A(n860), .B(n539), .CI(n814), .CO(n515), .S(n516) );
  CFA1X1 U424 ( .A(n839), .B(n761), .CI(n786), .CO(n517), .S(n518) );
  CFA1X1 U425 ( .A(n800), .B(n850), .CI(n773), .CO(n519), .S(n520) );
  CHA1X1 U426 ( .A(n750), .B(n827), .CO(n521), .S(n522) );
  CFA1X1 U427 ( .A(n528), .B(n526), .CI(n543), .CO(n523), .S(n524) );
  CFA1X1 U428 ( .A(n532), .B(n545), .CI(n530), .CO(n525), .S(n526) );
  CFA1X1 U429 ( .A(n534), .B(n547), .CI(n549), .CO(n527), .S(n528) );
  CFA1X1 U430 ( .A(n551), .B(n536), .CI(n538), .CO(n529), .S(n530) );
  CFA1X1 U431 ( .A(n555), .B(n553), .CI(n540), .CO(n531), .S(n532) );
  CFA1X1 U432 ( .A(n840), .B(n828), .CI(n851), .CO(n533), .S(n534) );
  CFA1X1 U433 ( .A(n815), .B(n774), .CI(n870), .CO(n535), .S(n536) );
  CFA1X1 U434 ( .A(n787), .B(n801), .CI(n861), .CO(n537), .S(n538) );
  CHA1X1 U435 ( .A(a[10]), .B(n762), .CO(n539), .S(n540) );
  CFA1X1 U436 ( .A(n546), .B(n544), .CI(n559), .CO(n541), .S(n542) );
  CFA1X1 U437 ( .A(n563), .B(n548), .CI(n561), .CO(n543), .S(n544) );
  CFA1X1 U438 ( .A(n554), .B(n550), .CI(n552), .CO(n545), .S(n546) );
  CFA1X1 U439 ( .A(n569), .B(n565), .CI(n567), .CO(n547), .S(n548) );
  CFA1X1 U440 ( .A(n841), .B(n556), .CI(n571), .CO(n549), .S(n550) );
  CFA1X1 U441 ( .A(n862), .B(n788), .CI(n816), .CO(n551), .S(n552) );
  CFA1X1 U442 ( .A(n871), .B(n829), .CI(n802), .CO(n553), .S(n554) );
  CHA1X1 U443 ( .A(n775), .B(n852), .CO(n555), .S(n556) );
  CFA1X1 U444 ( .A(n562), .B(n560), .CI(n575), .CO(n557), .S(n558) );
  CFA1X1 U445 ( .A(n579), .B(n564), .CI(n577), .CO(n559), .S(n560) );
  CFA1X1 U446 ( .A(n570), .B(n566), .CI(n568), .CO(n561), .S(n562) );
  CFA1X1 U447 ( .A(n572), .B(n581), .CI(n583), .CO(n563), .S(n564) );
  CFA1X1 U448 ( .A(n872), .B(n585), .CI(n853), .CO(n565), .S(n566) );
  CFA1X1 U449 ( .A(n817), .B(n803), .CI(n880), .CO(n567), .S(n568) );
  CHA1X1 U451 ( .A(n789), .B(n863), .CO(n571), .S(n572) );
  CFA1X1 U452 ( .A(n578), .B(n576), .CI(n589), .CO(n573), .S(n574) );
  CFA1X1 U453 ( .A(n593), .B(n591), .CI(n580), .CO(n575), .S(n576) );
  CFA1X1 U454 ( .A(n597), .B(n582), .CI(n584), .CO(n577), .S(n578) );
  CFA1X1 U455 ( .A(n599), .B(n595), .CI(n586), .CO(n579), .S(n580) );
  CFA1X1 U456 ( .A(n881), .B(n818), .CI(n843), .CO(n581), .S(n582) );
  CFA1X1 U457 ( .A(n873), .B(n864), .CI(n854), .CO(n583), .S(n584) );
  CHA1X1 U458 ( .A(n804), .B(n831), .CO(n585), .S(n586) );
  CFA1X1 U459 ( .A(n592), .B(n590), .CI(n603), .CO(n587), .S(n588) );
  CFA1X1 U460 ( .A(n596), .B(n605), .CI(n594), .CO(n589), .S(n590) );
  CFA1X1 U461 ( .A(n609), .B(n598), .CI(n607), .CO(n591), .S(n592) );
  CFA1X1 U462 ( .A(n882), .B(n600), .CI(n611), .CO(n593), .S(n594) );
  CFA1X1 U463 ( .A(n865), .B(n855), .CI(n889), .CO(n595), .S(n596) );
  CFA1X1 U464 ( .A(n844), .B(n832), .CI(n874), .CO(n597), .S(n598) );
  CHA1X1 U465 ( .A(a[8]), .B(n819), .CO(n599), .S(n600) );
  CFA1X1 U466 ( .A(n606), .B(n604), .CI(n615), .CO(n601), .S(n602) );
  CFA1X1 U467 ( .A(n610), .B(n617), .CI(n608), .CO(n603), .S(n604) );
  CFA1X1 U468 ( .A(n612), .B(n621), .CI(n619), .CO(n605), .S(n606) );
  CFA1X1 U469 ( .A(n866), .B(n623), .CI(n845), .CO(n607), .S(n608) );
  CFA1X1 U470 ( .A(n856), .B(n883), .CI(n890), .CO(n609), .S(n610) );
  CHA1X1 U471 ( .A(n875), .B(n833), .CO(n611), .S(n612) );
  CFA1X1 U472 ( .A(n627), .B(n616), .CI(n618), .CO(n613), .S(n614) );
  CFA1X1 U473 ( .A(n622), .B(n629), .CI(n620), .CO(n615), .S(n616) );
  CFA1X1 U474 ( .A(n633), .B(n631), .CI(n624), .CO(n617), .S(n618) );
  CFA1X1 U475 ( .A(n867), .B(n876), .CI(n897), .CO(n619), .S(n620) );
  CFA1X1 U476 ( .A(n846), .B(n857), .CI(n891), .CO(n621), .S(n622) );
  CFA1X1 U478 ( .A(n630), .B(n628), .CI(n637), .CO(n625), .S(n626) );
  CFA1X1 U479 ( .A(n641), .B(n632), .CI(n639), .CO(n627), .S(n628) );
  CFA1X1 U480 ( .A(n868), .B(n634), .CI(n643), .CO(n629), .S(n630) );
  CFA1X1 U481 ( .A(n858), .B(n898), .CI(n885), .CO(n631), .S(n632) );
  CHA1X1 U482 ( .A(n877), .B(n892), .CO(n633), .S(n634) );
  CFA1X1 U483 ( .A(n640), .B(n638), .CI(n647), .CO(n635), .S(n636) );
  CFA1X1 U484 ( .A(n644), .B(n642), .CI(n649), .CO(n637), .S(n638) );
  CFA1X1 U485 ( .A(n899), .B(n651), .CI(n904), .CO(n639), .S(n640) );
  CFA1X1 U486 ( .A(n886), .B(n878), .CI(n893), .CO(n641), .S(n642) );
  CHA1X1 U487 ( .A(a[6]), .B(n869), .CO(n643), .S(n644) );
  CFA1X1 U488 ( .A(n650), .B(n648), .CI(n655), .CO(n645), .S(n646) );
  CFA1X1 U489 ( .A(n652), .B(n657), .CI(n659), .CO(n647), .S(n648) );
  CFA1X1 U490 ( .A(n905), .B(n887), .CI(n900), .CO(n649), .S(n650) );
  CHA1X1 U491 ( .A(n879), .B(n894), .CO(n651), .S(n652) );
  CFA1X1 U492 ( .A(n663), .B(n656), .CI(n658), .CO(n653), .S(n654) );
  CFA1X1 U493 ( .A(n910), .B(n660), .CI(n665), .CO(n655), .S(n656) );
  CFA1X1 U494 ( .A(n888), .B(n895), .CI(n906), .CO(n657), .S(n658) );
  CFA1X1 U496 ( .A(n671), .B(n664), .CI(n669), .CO(n661), .S(n662) );
  CFA1X1 U497 ( .A(n911), .B(n666), .CI(n902), .CO(n663), .S(n664) );
  CHA1X1 U498 ( .A(n896), .B(n907), .CO(n665), .S(n666) );
  CFA1X1 U499 ( .A(n675), .B(n670), .CI(n672), .CO(n667), .S(n668) );
  CFA1X1 U500 ( .A(n912), .B(n908), .CI(n915), .CO(n669), .S(n670) );
  CHA1X1 U501 ( .A(a[4]), .B(n903), .CO(n671), .S(n672) );
  CFA1X1 U502 ( .A(n913), .B(n679), .CI(n676), .CO(n673), .S(n674) );
  CHA1X1 U503 ( .A(n916), .B(n909), .CO(n675), .S(n676) );
  CFA1X1 U504 ( .A(n919), .B(n681), .CI(n917), .CO(n677), .S(n678) );
  CHA1X1 U506 ( .A(n918), .B(n920), .CO(n681), .S(n682) );
  CHA1X1 U507 ( .A(a[2]), .B(n921), .CO(n683), .S(n684) );
  CIVX2 U796 ( .A(\b[0] ), .Z(n32) );
  CANR1X1 U797 ( .A(n227), .B(n219), .C(n220), .Z(n218) );
  CANR1XL U798 ( .A(n1031), .B(n159), .C(n154), .Z(n152) );
  CANR1XL U799 ( .A(n1032), .B(n197), .C(n192), .Z(n190) );
  COND1XL U800 ( .A(n166), .B(n160), .C(n161), .Z(n159) );
  CANR1X1 U801 ( .A(n146), .B(n1025), .C(n139), .Z(n133) );
  CENX1 U802 ( .A(n110), .B(n63), .Z(product[28]) );
  CIVX2 U803 ( .A(b[7]), .Z(n1043) );
  CIVX2 U804 ( .A(b[11]), .Z(n1046) );
  CIVX2 U805 ( .A(b[6]), .Z(n44) );
  CIVX1 U806 ( .A(b[3]), .Z(n1041) );
  COR2X1 U807 ( .A(n444), .B(n465), .Z(n1025) );
  COR2X1 U808 ( .A(n924), .B(a[1]), .Z(n1026) );
  CFA1XL U809 ( .A(a[11]), .B(n826), .CI(n785), .CO(n499), .S(n500) );
  CIVX1 U810 ( .A(b[14]), .Z(n949) );
  CENXL U811 ( .A(n103), .B(n62), .Z(product[29]) );
  CNR2XL U812 ( .A(n951), .B(n18), .Z(n763) );
  CIVX2 U813 ( .A(b[12]), .Z(n951) );
  CENXL U814 ( .A(n1027), .B(n89), .Z(product[31]) );
  CIVX2 U815 ( .A(b[16]), .Z(n16) );
  COND1X1 U816 ( .A(n206), .B(n189), .C(n190), .Z(n188) );
  CND2XL U817 ( .A(n196), .B(n1032), .Z(n189) );
  CIVX1 U818 ( .A(n141), .Z(n139) );
  CNR2XL U819 ( .A(n198), .B(n203), .Z(n196) );
  CIVX1 U820 ( .A(b[8]), .Z(n48) );
  CENX1 U821 ( .A(n122), .B(n65), .Z(product[26]) );
  CNR2XL U822 ( .A(n221), .B(n224), .Z(n219) );
  CND2XL U823 ( .A(n506), .B(n523), .Z(n161) );
  CND2IXL U824 ( .B(n111), .A(n112), .Z(n64) );
  CIVXL U825 ( .A(n132), .Z(n134) );
  CIVX1 U826 ( .A(n143), .Z(n258) );
  CNR2X1 U827 ( .A(n506), .B(n523), .Z(n160) );
  CANR1XL U828 ( .A(n1035), .B(n235), .C(n232), .Z(n230) );
  CNR2XL U829 ( .A(n44), .B(n48), .Z(n890) );
  CNR2XL U830 ( .A(n1044), .B(n20), .Z(n741) );
  CNR2XL U831 ( .A(n40), .B(n44), .Z(n905) );
  CNR2XL U832 ( .A(n1047), .B(n949), .Z(n820) );
  CNR2XL U833 ( .A(n1047), .B(n16), .Z(n791) );
  CNR2XL U834 ( .A(n1045), .B(n16), .Z(n795) );
  CIVX1 U835 ( .A(b[10]), .Z(n52) );
  CNR2X1 U836 ( .A(n1041), .B(n949), .Z(n830) );
  CANR1X1 U837 ( .A(n150), .B(n114), .C(n115), .Z(n59) );
  CNR2XL U838 ( .A(n116), .B(n132), .Z(n114) );
  CND2XL U839 ( .A(n1029), .B(n1030), .Z(n116) );
  COND1X1 U840 ( .A(n151), .B(n168), .C(n152), .Z(n150) );
  CND2XL U841 ( .A(n158), .B(n1031), .Z(n151) );
  CEOXL U842 ( .A(n70), .B(n162), .Z(product[21]) );
  CEOXL U843 ( .A(n68), .B(n149), .Z(product[23]) );
  CND2XL U844 ( .A(n258), .B(n144), .Z(n68) );
  CEOXL U845 ( .A(n69), .B(n157), .Z(product[22]) );
  CND2XL U846 ( .A(n1031), .B(n156), .Z(n69) );
  CND2XL U847 ( .A(n264), .B(n182), .Z(n74) );
  CND2XL U848 ( .A(n1032), .B(n194), .Z(n75) );
  CND2XL U849 ( .A(n261), .B(n166), .Z(n71) );
  CND2XL U850 ( .A(n1029), .B(n121), .Z(n65) );
  CND2XL U851 ( .A(n134), .B(n1030), .Z(n123) );
  CND2XL U852 ( .A(n348), .B(n373), .Z(n109) );
  CND2XL U853 ( .A(n294), .B(n321), .Z(n95) );
  CANR1X1 U854 ( .A(n207), .B(n215), .C(n208), .Z(n206) );
  CNR2XL U855 ( .A(n212), .B(n209), .Z(n207) );
  COND1X1 U856 ( .A(n216), .B(n218), .C(n217), .Z(n215) );
  CNR2XL U857 ( .A(n574), .B(n587), .Z(n181) );
  CNR2XL U858 ( .A(n466), .B(n485), .Z(n143) );
  CND2XL U859 ( .A(n269), .B(n213), .Z(n79) );
  CND2XL U860 ( .A(n270), .B(n217), .Z(n80) );
  CND2XL U861 ( .A(n267), .B(n204), .Z(n77) );
  CND2XL U862 ( .A(n1033), .B(n179), .Z(n73) );
  CND2XL U863 ( .A(n1033), .B(n264), .Z(n174) );
  CIVXL U864 ( .A(n203), .Z(n267) );
  CIVXL U865 ( .A(n204), .Z(n202) );
  CENX1 U866 ( .A(n279), .B(n293), .Z(n1027) );
  CND2XL U867 ( .A(n271), .B(n222), .Z(n81) );
  CND2XL U868 ( .A(n626), .B(n635), .Z(n210) );
  CND2XL U869 ( .A(n602), .B(n613), .Z(n199) );
  CND2XL U870 ( .A(n542), .B(n557), .Z(n172) );
  CND2XL U871 ( .A(n273), .B(n229), .Z(n83) );
  CEOXL U872 ( .A(n230), .B(n83), .Z(product[8]) );
  CND2XL U873 ( .A(n1035), .B(n234), .Z(n84) );
  CND2XL U874 ( .A(n272), .B(n225), .Z(n82) );
  COAN1XL U875 ( .A(n240), .B(n242), .C(n241), .Z(n1034) );
  CEOXL U876 ( .A(n1034), .B(n85), .Z(product[6]) );
  CND2XL U877 ( .A(n276), .B(n241), .Z(n86) );
  CEOXL U878 ( .A(n242), .B(n86), .Z(product[5]) );
  CND2XL U879 ( .A(n1028), .B(n246), .Z(n87) );
  CNR2XL U880 ( .A(n1048), .B(n40), .Z(n815) );
  CNR2XL U881 ( .A(n1048), .B(n36), .Z(n817) );
  CNR2XL U882 ( .A(n1040), .B(n23), .Z(n717) );
  CNR2XL U883 ( .A(n1040), .B(n1048), .Z(n816) );
  CNR2XL U884 ( .A(n1046), .B(n1048), .Z(n808) );
  CIVX1 U885 ( .A(b[5]), .Z(n1042) );
  CNR2XL U886 ( .A(n1042), .B(n18), .Z(n770) );
  CNR2XL U887 ( .A(n1042), .B(n22), .Z(n724) );
  COR2X1 U888 ( .A(n684), .B(n922), .Z(n1028) );
  CNR2XL U889 ( .A(n1043), .B(n951), .Z(n851) );
  CNR2XL U890 ( .A(n1042), .B(n949), .Z(n828) );
  CNR2XL U891 ( .A(n1043), .B(n21), .Z(n732) );
  CNR2XL U892 ( .A(n1040), .B(n25), .Z(n702) );
  CNR2XL U893 ( .A(n1041), .B(n48), .Z(n893) );
  CNR2XL U894 ( .A(n1043), .B(n19), .Z(n755) );
  CNR2XL U895 ( .A(n1042), .B(n21), .Z(n734) );
  CNR2XL U896 ( .A(n1048), .B(n44), .Z(n813) );
  CNR2XL U897 ( .A(n1043), .B(n1048), .Z(n812) );
  CNR2XL U898 ( .A(n1040), .B(n21), .Z(n736) );
  CNR2XL U899 ( .A(n1041), .B(n18), .Z(n772) );
  CNR2XL U900 ( .A(n1042), .B(n1044), .Z(n883) );
  CNR2XL U901 ( .A(n1048), .B(n52), .Z(n809) );
  CNR2XL U902 ( .A(n1041), .B(n20), .Z(n747) );
  CNR2XL U903 ( .A(n1040), .B(n22), .Z(n726) );
  CNR2XL U904 ( .A(n1042), .B(n48), .Z(n891) );
  CNR2XL U905 ( .A(n1048), .B(n951), .Z(n807) );
  CNR2XL U906 ( .A(n1040), .B(n26), .Z(n696) );
  CNR2XL U907 ( .A(n1041), .B(n16), .Z(n801) );
  CNR2XL U908 ( .A(n1041), .B(n17), .Z(n786) );
  CNR2XL U909 ( .A(n1043), .B(n1047), .Z(n839) );
  CNR2XL U910 ( .A(n1041), .B(n1046), .Z(n866) );
  CNR2XL U911 ( .A(n1038), .B(n1047), .Z(n845) );
  CNR2XL U912 ( .A(n1041), .B(n52), .Z(n876) );
  CNR2XL U913 ( .A(n1043), .B(n44), .Z(n897) );
  CNR2XL U914 ( .A(n1041), .B(n1043), .Z(n900) );
  CNR2XL U915 ( .A(n1042), .B(n23), .Z(n715) );
  CNR2XL U916 ( .A(n1043), .B(n40), .Z(n899) );
  CNR2XL U917 ( .A(n1042), .B(n44), .Z(n904) );
  CNR2XL U918 ( .A(n1041), .B(n19), .Z(n759) );
  CNR2XL U919 ( .A(n1042), .B(n17), .Z(n784) );
  CNR2XL U920 ( .A(n1040), .B(n24), .Z(n709) );
  CNR2XL U921 ( .A(n1042), .B(n1046), .Z(n864) );
  CNR2XL U922 ( .A(n1042), .B(n20), .Z(n745) );
  CNR2XL U923 ( .A(n1042), .B(n19), .Z(n757) );
  CNR2XL U924 ( .A(n1047), .B(n1048), .Z(n806) );
  CNR2XL U925 ( .A(n1042), .B(n24), .Z(n707) );
  CNR2XL U926 ( .A(n1041), .B(n951), .Z(n855) );
  CNR2XL U927 ( .A(n1042), .B(n1048), .Z(n814) );
  CNR2XL U928 ( .A(n1041), .B(n1044), .Z(n885) );
  CNR2XL U929 ( .A(n1042), .B(n1043), .Z(n898) );
  CNR2XL U930 ( .A(n1042), .B(n951), .Z(n853) );
  CNR2XL U931 ( .A(n1044), .B(n1048), .Z(n810) );
  CNR2XL U932 ( .A(n1048), .B(n949), .Z(n805) );
  CNR2XL U933 ( .A(n1041), .B(n1047), .Z(n843) );
  CNR2XL U934 ( .A(n1042), .B(n52), .Z(n874) );
  CNR2XL U935 ( .A(n1043), .B(n20), .Z(n743) );
  CNR2XL U936 ( .A(n1043), .B(n22), .Z(n722) );
  CNR2XL U937 ( .A(n1042), .B(n25), .Z(n700) );
  CND2XL U938 ( .A(n678), .B(n680), .Z(n237) );
  CNR2XL U939 ( .A(n1040), .B(n36), .Z(n919) );
  CNR2XL U940 ( .A(n1038), .B(n40), .Z(n917) );
  CNR2XL U941 ( .A(n1041), .B(n27), .Z(n691) );
  CEOXL U942 ( .A(n1036), .B(n250), .Z(product[3]) );
  CIVX1 U943 ( .A(b[2]), .Z(n36) );
  CIVX1 U944 ( .A(b[4]), .Z(n40) );
  CNR2XL U945 ( .A(n1047), .B(n40), .Z(n842) );
  CIVXL U946 ( .A(b[17]), .Z(n17) );
  CIVXL U947 ( .A(b[18]), .Z(n18) );
  CNR2XL U948 ( .A(n1045), .B(n40), .Z(n884) );
  CIVXL U949 ( .A(b[20]), .Z(n20) );
  CIVXL U950 ( .A(b[21]), .Z(n21) );
  CIVXL U951 ( .A(b[22]), .Z(n22) );
  CNR2XL U952 ( .A(n1046), .B(n32), .Z(n869) );
  CNR2XL U953 ( .A(n23), .B(n32), .Z(n720) );
  CNR2XL U954 ( .A(n1043), .B(n949), .Z(n826) );
  CNR2XL U955 ( .A(n17), .B(n40), .Z(n785) );
  CNR2XL U956 ( .A(n1042), .B(n32), .Z(n914) );
  CNR2XL U957 ( .A(n1043), .B(n32), .Z(n903) );
  CNR2XL U958 ( .A(n19), .B(n32), .Z(n762) );
  CNR2XL U959 ( .A(n1048), .B(n32), .Z(n819) );
  CNR2XL U960 ( .A(n27), .B(n32), .Z(n694) );
  CIVXL U961 ( .A(b[28]), .Z(n28) );
  CNR2XL U962 ( .A(n32), .B(n30), .Z(n685) );
  CAN2XL U963 ( .A(n1026), .B(n250), .Z(product[2]) );
  CND2X1 U964 ( .A(n106), .B(n99), .Z(n97) );
  CND2X1 U965 ( .A(n92), .B(n106), .Z(n90) );
  COND1XL U966 ( .A(n112), .B(n108), .C(n109), .Z(n107) );
  CNR2X1 U967 ( .A(n108), .B(n111), .Z(n106) );
  CANR1XL U968 ( .A(n99), .B(n107), .C(n100), .Z(n98) );
  CANR1XL U969 ( .A(n107), .B(n92), .C(n93), .Z(n91) );
  COND1XL U970 ( .A(n102), .B(n94), .C(n95), .Z(n93) );
  CANR1XL U971 ( .A(n128), .B(n1029), .C(n119), .Z(n117) );
  CND2X1 U972 ( .A(n253), .B(n109), .Z(n63) );
  COND1XL U973 ( .A(n111), .B(n59), .C(n112), .Z(n110) );
  CND2X1 U974 ( .A(n99), .B(n102), .Z(n62) );
  COND1XL U975 ( .A(n104), .B(n59), .C(n105), .Z(n103) );
  CENX1 U976 ( .A(n96), .B(n61), .Z(product[30]) );
  CND2X1 U977 ( .A(n251), .B(n95), .Z(n61) );
  COND1XL U978 ( .A(n97), .B(n59), .C(n98), .Z(n96) );
  CNR2X1 U979 ( .A(n94), .B(n101), .Z(n92) );
  COND1XL U980 ( .A(n133), .B(n116), .C(n117), .Z(n115) );
  CNR2X1 U981 ( .A(n374), .B(n397), .Z(n111) );
  CNR2X1 U982 ( .A(n348), .B(n373), .Z(n108) );
  CNR2X1 U983 ( .A(n294), .B(n321), .Z(n94) );
  CANR1XL U984 ( .A(n1030), .B(n135), .C(n128), .Z(n124) );
  CNR2X1 U985 ( .A(n322), .B(n347), .Z(n101) );
  CENX1 U986 ( .A(n131), .B(n66), .Z(product[25]) );
  CND2X1 U987 ( .A(n1030), .B(n130), .Z(n66) );
  COND1XL U988 ( .A(n132), .B(n149), .C(n133), .Z(n131) );
  CENX1 U989 ( .A(n142), .B(n67), .Z(product[24]) );
  CND2X1 U990 ( .A(n1025), .B(n141), .Z(n67) );
  COND1XL U991 ( .A(n143), .B(n149), .C(n144), .Z(n142) );
  COND1XL U992 ( .A(n123), .B(n149), .C(n124), .Z(n122) );
  CENX1 U993 ( .A(n167), .B(n71), .Z(product[20]) );
  CNR2X1 U994 ( .A(n160), .B(n165), .Z(n158) );
  CANR1XL U995 ( .A(n158), .B(n167), .C(n159), .Z(n157) );
  CEOX1 U996 ( .A(n74), .B(n187), .Z(product[17]) );
  CEOX1 U997 ( .A(n75), .B(n195), .Z(product[16]) );
  CANR1XL U998 ( .A(n196), .B(n205), .C(n197), .Z(n195) );
  CND2X1 U999 ( .A(n260), .B(n161), .Z(n70) );
  CANR1XL U1000 ( .A(n261), .B(n167), .C(n164), .Z(n162) );
  COR2X1 U1001 ( .A(n398), .B(n421), .Z(n1029) );
  CND2X1 U1002 ( .A(n322), .B(n347), .Z(n102) );
  CND2X1 U1003 ( .A(n1025), .B(n258), .Z(n132) );
  CND2X1 U1004 ( .A(n374), .B(n397), .Z(n112) );
  CND2X1 U1005 ( .A(n398), .B(n421), .Z(n121) );
  COND1XL U1006 ( .A(n213), .B(n209), .C(n210), .Z(n208) );
  CNR2X1 U1007 ( .A(n174), .B(n171), .Z(n169) );
  COND1XL U1008 ( .A(n171), .B(n175), .C(n172), .Z(n170) );
  CANR1XL U1009 ( .A(n184), .B(n1033), .C(n177), .Z(n175) );
  COND1XL U1010 ( .A(n204), .B(n198), .C(n199), .Z(n197) );
  CNR2X1 U1011 ( .A(n524), .B(n541), .Z(n165) );
  COR2X1 U1012 ( .A(n422), .B(n443), .Z(n1030) );
  CENX1 U1013 ( .A(n211), .B(n78), .Z(product[13]) );
  CND2X1 U1014 ( .A(n268), .B(n210), .Z(n78) );
  COND1XL U1015 ( .A(n212), .B(n214), .C(n213), .Z(n211) );
  CENX1 U1016 ( .A(n205), .B(n77), .Z(product[14]) );
  CENX1 U1017 ( .A(n180), .B(n73), .Z(product[18]) );
  COND1XL U1018 ( .A(n181), .B(n187), .C(n182), .Z(n180) );
  CND2X1 U1019 ( .A(n262), .B(n172), .Z(n72) );
  COND1XL U1020 ( .A(n174), .B(n187), .C(n175), .Z(n173) );
  CEOX1 U1021 ( .A(n76), .B(n200), .Z(product[15]) );
  CND2X1 U1022 ( .A(n266), .B(n199), .Z(n76) );
  CANR1XL U1023 ( .A(n267), .B(n205), .C(n202), .Z(n200) );
  CEOX1 U1024 ( .A(n80), .B(n218), .Z(product[11]) );
  CEOX1 U1025 ( .A(n79), .B(n214), .Z(product[12]) );
  COR2X1 U1026 ( .A(n486), .B(n505), .Z(n1031) );
  COR2X1 U1027 ( .A(n588), .B(n601), .Z(n1032) );
  CND2X1 U1028 ( .A(n466), .B(n485), .Z(n144) );
  CND2X1 U1029 ( .A(n574), .B(n587), .Z(n182) );
  CND2X1 U1030 ( .A(n524), .B(n541), .Z(n166) );
  CND2X1 U1031 ( .A(n422), .B(n443), .Z(n130) );
  CND2X1 U1032 ( .A(n444), .B(n465), .Z(n141) );
  CND2X1 U1033 ( .A(n486), .B(n505), .Z(n156) );
  CND2X1 U1034 ( .A(n588), .B(n601), .Z(n194) );
  COND1XL U1035 ( .A(n225), .B(n221), .C(n222), .Z(n220) );
  COND1XL U1036 ( .A(n230), .B(n228), .C(n229), .Z(n227) );
  CNR2X1 U1037 ( .A(n542), .B(n557), .Z(n171) );
  CNR2X1 U1038 ( .A(n626), .B(n635), .Z(n209) );
  CNR2X1 U1039 ( .A(n636), .B(n645), .Z(n212) );
  CNR2X1 U1040 ( .A(n602), .B(n613), .Z(n198) );
  CNR2X1 U1041 ( .A(n614), .B(n625), .Z(n203) );
  CENX1 U1042 ( .A(n81), .B(n223), .Z(product[10]) );
  COND1XL U1043 ( .A(n224), .B(n226), .C(n225), .Z(n223) );
  CNR2X1 U1044 ( .A(n646), .B(n653), .Z(n216) );
  COND1XL U1045 ( .A(n90), .B(n59), .C(n91), .Z(n89) );
  COR2X1 U1046 ( .A(n558), .B(n573), .Z(n1033) );
  CND2X1 U1047 ( .A(n614), .B(n625), .Z(n204) );
  CND2X1 U1048 ( .A(n636), .B(n645), .Z(n213) );
  CND2X1 U1049 ( .A(n558), .B(n573), .Z(n179) );
  CND2X1 U1050 ( .A(n646), .B(n653), .Z(n217) );
  CENX1 U1051 ( .A(n235), .B(n84), .Z(product[7]) );
  CEOX1 U1052 ( .A(n226), .B(n82), .Z(product[9]) );
  CANR1XL U1053 ( .A(n247), .B(n1028), .C(n244), .Z(n242) );
  COND1XL U1054 ( .A(n1034), .B(n236), .C(n237), .Z(n235) );
  CNR2X1 U1055 ( .A(n662), .B(n667), .Z(n224) );
  CNR2X1 U1056 ( .A(n654), .B(n661), .Z(n221) );
  CNR2X1 U1057 ( .A(n668), .B(n673), .Z(n228) );
  CNR2X1 U1058 ( .A(n1042), .B(n1047), .Z(n841) );
  CND2X1 U1059 ( .A(n662), .B(n667), .Z(n225) );
  CND2X1 U1060 ( .A(n674), .B(n677), .Z(n234) );
  CND2X1 U1061 ( .A(n654), .B(n661), .Z(n222) );
  CND2X1 U1062 ( .A(n668), .B(n673), .Z(n229) );
  COR2X1 U1063 ( .A(n674), .B(n677), .Z(n1035) );
  CND2X1 U1064 ( .A(n275), .B(n237), .Z(n85) );
  CNR2X1 U1065 ( .A(n25), .B(n32), .Z(n705) );
  CNR2X1 U1066 ( .A(n1043), .B(n36), .Z(n901) );
  CNR2X1 U1067 ( .A(n40), .B(n949), .Z(n829) );
  CNR2X1 U1068 ( .A(n36), .B(n16), .Z(n802) );
  CNR2X1 U1069 ( .A(n48), .B(n52), .Z(n871) );
  CNR2X1 U1070 ( .A(n951), .B(n52), .Z(n848) );
  CNR2X1 U1071 ( .A(n32), .B(n22), .Z(n729) );
  CNR2X1 U1072 ( .A(n40), .B(n18), .Z(n771) );
  CNR2X1 U1073 ( .A(n1047), .B(n32), .Z(n846) );
  CNR2X1 U1074 ( .A(n1047), .B(n36), .Z(n844) );
  CNR2X1 U1075 ( .A(n17), .B(n951), .Z(n777) );
  CNR2X1 U1076 ( .A(n21), .B(n48), .Z(n731) );
  CNR2X1 U1077 ( .A(n25), .B(n40), .Z(n701) );
  CNR2X1 U1078 ( .A(n1046), .B(n18), .Z(n764) );
  CNR2X1 U1079 ( .A(n48), .B(n951), .Z(n850) );
  CNR2X1 U1080 ( .A(n40), .B(n16), .Z(n800) );
  CNR2X1 U1081 ( .A(n36), .B(n18), .Z(n773) );
  CNR2X1 U1082 ( .A(n36), .B(n24), .Z(n710) );
  CNR2X1 U1083 ( .A(n32), .B(n26), .Z(n699) );
  CNR2X1 U1084 ( .A(n48), .B(n18), .Z(n767) );
  CNR2X1 U1085 ( .A(n19), .B(n48), .Z(n754) );
  CNR2X1 U1086 ( .A(n1047), .B(n44), .Z(n840) );
  CNR2X1 U1087 ( .A(n1043), .B(n1046), .Z(n862) );
  CNR2X1 U1088 ( .A(n17), .B(n52), .Z(n779) );
  CNR2X1 U1089 ( .A(n23), .B(n40), .Z(n716) );
  CNR2X1 U1090 ( .A(n1046), .B(n16), .Z(n793) );
  CNR2X1 U1091 ( .A(n36), .B(n951), .Z(n856) );
  CNR2X1 U1092 ( .A(n21), .B(n36), .Z(n737) );
  CNR2X1 U1093 ( .A(n1048), .B(n48), .Z(n811) );
  CNR2X1 U1094 ( .A(n1045), .B(n949), .Z(n824) );
  CNR2X1 U1095 ( .A(n1043), .B(n16), .Z(n797) );
  CNR2X1 U1096 ( .A(n1044), .B(n19), .Z(n753) );
  CNR2X1 U1097 ( .A(n1045), .B(n36), .Z(n886) );
  CNR2X1 U1098 ( .A(n19), .B(n44), .Z(n756) );
  CNR2X1 U1099 ( .A(n1047), .B(n951), .Z(n834) );
  CNR2X1 U1100 ( .A(n682), .B(n683), .Z(n240) );
  CNR2X1 U1101 ( .A(n678), .B(n680), .Z(n236) );
  CNR2X1 U1102 ( .A(n1042), .B(n16), .Z(n799) );
  CNR2X1 U1103 ( .A(n1047), .B(n48), .Z(n838) );
  CNR2X1 U1104 ( .A(n19), .B(n36), .Z(n760) );
  CNR2X1 U1105 ( .A(n21), .B(n44), .Z(n733) );
  CNR2X1 U1106 ( .A(n25), .B(n36), .Z(n703) );
  CNR2X1 U1107 ( .A(n1043), .B(n17), .Z(n782) );
  CNR2X1 U1108 ( .A(n17), .B(n36), .Z(n787) );
  CNR2X1 U1109 ( .A(n1046), .B(n48), .Z(n861) );
  CNR2X1 U1110 ( .A(n1044), .B(n48), .Z(n880) );
  CNR2X1 U1111 ( .A(n23), .B(n36), .Z(n718) );
  CNR2X1 U1112 ( .A(n17), .B(n48), .Z(n781) );
  CNR2X1 U1113 ( .A(n1046), .B(n949), .Z(n822) );
  CNR2X1 U1114 ( .A(n1046), .B(n36), .Z(n867) );
  CNR2X1 U1115 ( .A(n1043), .B(n18), .Z(n768) );
  CNR2X1 U1116 ( .A(n52), .B(n16), .Z(n794) );
  CNR2X1 U1117 ( .A(n40), .B(n22), .Z(n725) );
  CNR2X1 U1118 ( .A(n1046), .B(n17), .Z(n778) );
  CNR2X1 U1119 ( .A(n1047), .B(n52), .Z(n836) );
  CNR2X1 U1120 ( .A(n19), .B(n40), .Z(n758) );
  CNR2X1 U1121 ( .A(n44), .B(n22), .Z(n723) );
  CNR2X1 U1122 ( .A(n32), .B(n28), .Z(n690) );
  CNR2X1 U1123 ( .A(n52), .B(n18), .Z(n765) );
  CNR2X1 U1124 ( .A(n1046), .B(n44), .Z(n863) );
  CNR2X1 U1125 ( .A(n17), .B(n32), .Z(n789) );
  CNR2X1 U1126 ( .A(n23), .B(n44), .Z(n714) );
  CNR2X1 U1127 ( .A(n29), .B(n32), .Z(n687) );
  CNR2X1 U1128 ( .A(n40), .B(n52), .Z(n875) );
  CNR2X1 U1129 ( .A(n32), .B(n949), .Z(n833) );
  CNR2X1 U1130 ( .A(n44), .B(n20), .Z(n744) );
  CNR2X1 U1131 ( .A(n951), .B(n949), .Z(n821) );
  CNR2X1 U1132 ( .A(n44), .B(n52), .Z(n873) );
  CNR2X1 U1133 ( .A(n40), .B(n951), .Z(n854) );
  CNR2X1 U1134 ( .A(n1044), .B(n44), .Z(n882) );
  CNR2X1 U1135 ( .A(n1045), .B(n32), .Z(n888) );
  CNR2X1 U1136 ( .A(n1041), .B(n44), .Z(n906) );
  CNR2X1 U1137 ( .A(n951), .B(n16), .Z(n792) );
  CNR2X1 U1138 ( .A(n36), .B(n26), .Z(n697) );
  CNR2X1 U1139 ( .A(n19), .B(n52), .Z(n752) );
  CNR2X1 U1140 ( .A(n32), .B(n44), .Z(n909) );
  CNR2X1 U1141 ( .A(n36), .B(n40), .Z(n916) );
  CNR2X1 U1142 ( .A(n36), .B(n949), .Z(n831) );
  CNR2X1 U1143 ( .A(n32), .B(n16), .Z(n804) );
  CNR2X1 U1144 ( .A(n36), .B(n48), .Z(n894) );
  CNR2X1 U1145 ( .A(n32), .B(n52), .Z(n879) );
  CNR2X1 U1146 ( .A(n44), .B(n949), .Z(n827) );
  CNR2X1 U1147 ( .A(n32), .B(n20), .Z(n750) );
  CNR2X1 U1148 ( .A(n44), .B(n16), .Z(n798) );
  CNR2X1 U1149 ( .A(n1045), .B(n1047), .Z(n837) );
  CNR2X1 U1150 ( .A(n1045), .B(n52), .Z(n870) );
  CNR2X1 U1151 ( .A(n1046), .B(n40), .Z(n865) );
  CNR2X1 U1152 ( .A(n1043), .B(n48), .Z(n889) );
  CNR2X1 U1153 ( .A(n32), .B(n951), .Z(n858) );
  CNR2X1 U1154 ( .A(n1043), .B(n52), .Z(n872) );
  CNR2X1 U1155 ( .A(n21), .B(n40), .Z(n735) );
  CNR2X1 U1156 ( .A(n1044), .B(n18), .Z(n766) );
  CNR2X1 U1157 ( .A(n17), .B(n44), .Z(n783) );
  CNR2X1 U1158 ( .A(n1046), .B(n951), .Z(n847) );
  CNR2X1 U1159 ( .A(n1045), .B(n17), .Z(n780) );
  CNR2X1 U1160 ( .A(n1045), .B(n1046), .Z(n860) );
  CNR2X1 U1161 ( .A(n949), .B(n52), .Z(n823) );
  CNR2X1 U1162 ( .A(n48), .B(n16), .Z(n796) );
  CNR2X1 U1163 ( .A(n44), .B(n18), .Z(n769) );
  CNR2X1 U1164 ( .A(n48), .B(n20), .Z(n742) );
  CNR2X1 U1165 ( .A(n40), .B(n24), .Z(n708) );
  CNR2X1 U1166 ( .A(n32), .B(n40), .Z(n918) );
  CNR2X1 U1167 ( .A(n36), .B(n20), .Z(n748) );
  CNR2X1 U1168 ( .A(n48), .B(n949), .Z(n825) );
  CNR2X1 U1169 ( .A(n1046), .B(n52), .Z(n859) );
  CNR2X1 U1170 ( .A(n1045), .B(n951), .Z(n849) );
  CNR2X1 U1171 ( .A(n1041), .B(n1042), .Z(n911) );
  CNR2X1 U1172 ( .A(n1043), .B(n1044), .Z(n881) );
  CNR2X1 U1173 ( .A(n36), .B(n22), .Z(n727) );
  CNR2X1 U1174 ( .A(n1046), .B(n1047), .Z(n835) );
  CNR2X1 U1175 ( .A(n1042), .B(n40), .Z(n910) );
  CNR2X1 U1176 ( .A(n27), .B(n36), .Z(n692) );
  CNR2X1 U1177 ( .A(n1042), .B(n36), .Z(n912) );
  CNR2X1 U1178 ( .A(n1041), .B(n40), .Z(n915) );
  CNR2X1 U1179 ( .A(n21), .B(n32), .Z(n739) );
  CNR2X1 U1180 ( .A(n36), .B(n52), .Z(n877) );
  CNR2X1 U1181 ( .A(n40), .B(n48), .Z(n892) );
  CNR2X1 U1182 ( .A(n44), .B(n951), .Z(n852) );
  CNR2X1 U1183 ( .A(n32), .B(n18), .Z(n775) );
  CNR2X1 U1184 ( .A(n36), .B(n44), .Z(n907) );
  CNR2X1 U1185 ( .A(n32), .B(n48), .Z(n896) );
  CNR2X1 U1186 ( .A(n40), .B(n20), .Z(n746) );
  CNR2X1 U1187 ( .A(n32), .B(n24), .Z(n712) );
  CNR2X1 U1188 ( .A(n1047), .B(n17), .Z(n776) );
  CEOX1 U1189 ( .A(n685), .B(n688), .Z(n292) );
  CNR2X1 U1190 ( .A(n1045), .B(n21), .Z(n730) );
  CNR2X1 U1191 ( .A(n1043), .B(n23), .Z(n713) );
  CNR2X1 U1192 ( .A(n1046), .B(n19), .Z(n751) );
  CNR2X1 U1193 ( .A(n44), .B(n24), .Z(n706) );
  CNR2X1 U1194 ( .A(n40), .B(n26), .Z(n695) );
  CNR2X1 U1195 ( .A(n48), .B(n22), .Z(n721) );
  CNR2X1 U1196 ( .A(n949), .B(n16), .Z(n790) );
  CNR2X1 U1197 ( .A(n52), .B(n20), .Z(n740) );
  CND2X1 U1198 ( .A(n682), .B(n683), .Z(n241) );
  COR2X1 U1199 ( .A(n32), .B(n36), .Z(n1036) );
  CNR2X1 U1200 ( .A(n36), .B(n28), .Z(n688) );
  CNR2X1 U1201 ( .A(n1040), .B(n32), .Z(n921) );
  CEOXL U1202 ( .A(n64), .B(n59), .Z(product[27]) );
  CIVX1 U1203 ( .A(b[19]), .Z(n19) );
  CNR2X1 U1204 ( .A(n250), .B(n1036), .Z(n247) );
  CNR2X1 U1205 ( .A(n1038), .B(n32), .Z(n924) );
  CNR2XL U1206 ( .A(n1038), .B(n1048), .Z(n818) );
  CNR2X1 U1207 ( .A(n1038), .B(n949), .Z(n832) );
  CNR2X1 U1208 ( .A(n1038), .B(n951), .Z(n857) );
  CNR2XL U1209 ( .A(n1038), .B(n1046), .Z(n868) );
  CNR2X1 U1210 ( .A(n1038), .B(n52), .Z(n878) );
  CNR2XL U1211 ( .A(n1038), .B(n1044), .Z(n887) );
  CNR2X1 U1212 ( .A(n1039), .B(n48), .Z(n895) );
  CNR2XL U1213 ( .A(n1038), .B(n1043), .Z(n902) );
  CNR2X1 U1214 ( .A(n1038), .B(n44), .Z(n908) );
  CNR2X1 U1215 ( .A(n1038), .B(n1042), .Z(n913) );
  CNR2X1 U1216 ( .A(n1038), .B(n1040), .Z(n920) );
  CNR2X1 U1217 ( .A(n1039), .B(n36), .Z(n922) );
  CNR2X1 U1218 ( .A(n1038), .B(n16), .Z(n803) );
  CNR2X1 U1219 ( .A(n1039), .B(n17), .Z(n788) );
  CNR2X1 U1220 ( .A(n1039), .B(n18), .Z(n774) );
  CNR2X1 U1221 ( .A(n1039), .B(n19), .Z(n761) );
  CNR2X1 U1222 ( .A(n1039), .B(n20), .Z(n749) );
  CNR2X1 U1223 ( .A(n1039), .B(n21), .Z(n738) );
  CNR2X1 U1224 ( .A(n1039), .B(n22), .Z(n728) );
  CNR2X1 U1225 ( .A(n1039), .B(n23), .Z(n719) );
  CNR2X1 U1226 ( .A(n1039), .B(n24), .Z(n711) );
  CNR2X1 U1227 ( .A(n1039), .B(n25), .Z(n704) );
  CNR2X1 U1228 ( .A(n1038), .B(n26), .Z(n698) );
  CNR2X1 U1229 ( .A(n1039), .B(n27), .Z(n693) );
  CNR2X1 U1230 ( .A(n1039), .B(n28), .Z(n689) );
  CNR2X1 U1231 ( .A(n1039), .B(n29), .Z(n686) );
  CENX1 U1232 ( .A(n87), .B(n247), .Z(product[4]) );
  CND2X1 U1233 ( .A(n684), .B(n922), .Z(n246) );
  CHA1XL U1234 ( .A(a[7]), .B(n884), .CO(n623), .S(n624) );
  CND2XL U1235 ( .A(n924), .B(a[1]), .Z(n250) );
  CIVX1 U1236 ( .A(b[13]), .Z(n1047) );
  CHA1XL U1237 ( .A(n705), .B(a[13]), .CO(n419), .S(n420) );
  CHA1XL U1238 ( .A(a[3]), .B(n914), .CO(n679), .S(n680) );
  CHA1XL U1239 ( .A(a[5]), .B(n901), .CO(n659), .S(n660) );
  CFA1XL U1240 ( .A(a[9]), .B(n830), .CI(n842), .CO(n569), .S(n570) );
  CENX1 U1241 ( .A(n173), .B(n72), .Z(product[19]) );
  CIVXL U1242 ( .A(b[1]), .Z(n1038) );
  CIVXL U1243 ( .A(b[1]), .Z(n1039) );
  CIVXL U1244 ( .A(b[3]), .Z(n1040) );
  CIVXL U1245 ( .A(b[9]), .Z(n1044) );
  CIVXL U1246 ( .A(b[9]), .Z(n1045) );
  CIVXL U1247 ( .A(b[15]), .Z(n1048) );
  CIVX2 U1248 ( .A(b[30]), .Z(n30) );
  CIVX2 U1249 ( .A(b[29]), .Z(n29) );
  CIVX2 U1250 ( .A(n240), .Z(n276) );
  CIVX2 U1251 ( .A(n236), .Z(n275) );
  CIVX2 U1252 ( .A(n228), .Z(n273) );
  CIVX2 U1253 ( .A(n224), .Z(n272) );
  CIVX2 U1254 ( .A(n221), .Z(n271) );
  CIVX2 U1255 ( .A(n216), .Z(n270) );
  CIVX2 U1256 ( .A(b[27]), .Z(n27) );
  CIVX2 U1257 ( .A(n212), .Z(n269) );
  CIVX2 U1258 ( .A(n209), .Z(n268) );
  CIVX2 U1259 ( .A(n198), .Z(n266) );
  CIVX2 U1260 ( .A(n171), .Z(n262) );
  CIVX2 U1261 ( .A(n160), .Z(n260) );
  CIVX2 U1262 ( .A(b[26]), .Z(n26) );
  CIVX2 U1263 ( .A(n108), .Z(n253) );
  CIVX2 U1264 ( .A(n101), .Z(n99) );
  CIVX2 U1265 ( .A(n94), .Z(n251) );
  CIVX2 U1266 ( .A(b[25]), .Z(n25) );
  CIVX2 U1267 ( .A(n246), .Z(n244) );
  CIVX2 U1268 ( .A(b[24]), .Z(n24) );
  CIVX2 U1269 ( .A(n234), .Z(n232) );
  CIVX2 U1270 ( .A(b[23]), .Z(n23) );
  CIVX2 U1271 ( .A(n227), .Z(n226) );
  CIVX2 U1272 ( .A(n215), .Z(n214) );
  CIVX2 U1273 ( .A(n206), .Z(n205) );
  CIVX2 U1274 ( .A(n194), .Z(n192) );
  CIVX2 U1275 ( .A(n188), .Z(n187) );
  CIVX2 U1276 ( .A(n182), .Z(n184) );
  CIVX2 U1277 ( .A(n181), .Z(n264) );
  CIVX2 U1278 ( .A(n179), .Z(n177) );
  CIVX2 U1279 ( .A(n168), .Z(n167) );
  CIVX2 U1280 ( .A(n166), .Z(n164) );
  CIVX2 U1281 ( .A(n165), .Z(n261) );
  CIVX2 U1282 ( .A(n156), .Z(n154) );
  CIVX2 U1283 ( .A(n150), .Z(n149) );
  CIVX2 U1284 ( .A(n144), .Z(n146) );
  CIVX2 U1285 ( .A(n133), .Z(n135) );
  CIVX2 U1286 ( .A(n130), .Z(n128) );
  CIVX2 U1287 ( .A(n121), .Z(n119) );
  CIVX2 U1288 ( .A(n107), .Z(n105) );
  CIVX2 U1289 ( .A(n106), .Z(n104) );
  CIVX2 U1290 ( .A(n102), .Z(n100) );
endmodule


module calc ( clk, rst, A, B, C, pushA, stopA, pushB, stopB, pushC, stopC, Z, 
        pushZ );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  output [31:0] Z;
  input clk, rst, pushA, pushB, pushC;
  output stopA, stopB, stopC, pushZ;
  wire   all_in, all_in1, all_in2, all_in3, all_in4, all_in5, all_in6, all_in7,
         N6, n13, n14, n15, n16, n18, n20, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926;
  wire   [31:0] res_temp;
  wire   [31:0] captA;
  wire   [31:0] captB;
  wire   [31:0] captC;
  wire   [31:0] f01;
  wire   [31:0] f02;
  wire   [31:0] f03;
  wire   [31:0] f11;
  wire   [31:0] f12;
  wire   [31:0] f13;
  wire   [31:0] f14;
  wire   [31:0] f15;
  wire   [31:0] f16;
  wire   [31:0] f17;
  wire   [31:0] f21;
  wire   [31:0] f22;
  wire   [31:0] f23;
  wire   [31:0] f24;
  wire   [31:0] f25;
  wire   [31:0] f26;
  wire   [31:0] f27;
  wire   [31:0] f30;
  wire   [31:0] f31;
  wire   [31:0] f32;
  wire   [31:0] f33;
  wire   [31:0] f34;
  wire   [31:0] f41;
  wire   [31:0] f42;
  wire   [31:0] f43;
  wire   [31:0] f51;
  wire   [31:0] f52;
  wire   [31:0] res_d;
  wire   [2:0] seen_d;
  wire   [31:0] s12;
  wire   [31:0] s14;
  wire   [31:0] s15;
  wire   [31:0] s16;
  wire   [31:0] s17;
  wire   [31:0] s22;
  wire   [31:0] s23;
  wire   [31:0] s24;
  wire   [31:0] s26;
  wire   [31:0] s27;
  wire   [31:0] s31;
  wire   [31:0] s32;
  wire   [31:0] s33;
  wire   [31:0] s41;
  wire   [31:0] s43;
  wire   [31:0] s51;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, 
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        SYNOPSYS_UNCONNECTED__174, SYNOPSYS_UNCONNECTED__175, 
        SYNOPSYS_UNCONNECTED__176, SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, 
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        SYNOPSYS_UNCONNECTED__184, SYNOPSYS_UNCONNECTED__185, 
        SYNOPSYS_UNCONNECTED__186, SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, 
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, 
        SYNOPSYS_UNCONNECTED__202, SYNOPSYS_UNCONNECTED__203, 
        SYNOPSYS_UNCONNECTED__204, SYNOPSYS_UNCONNECTED__205, 
        SYNOPSYS_UNCONNECTED__206, SYNOPSYS_UNCONNECTED__207, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, 
        SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213, 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        SYNOPSYS_UNCONNECTED__216, SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, 
        SYNOPSYS_UNCONNECTED__222, SYNOPSYS_UNCONNECTED__223, 
        SYNOPSYS_UNCONNECTED__224, SYNOPSYS_UNCONNECTED__225, 
        SYNOPSYS_UNCONNECTED__226, SYNOPSYS_UNCONNECTED__227, 
        SYNOPSYS_UNCONNECTED__228, SYNOPSYS_UNCONNECTED__229, 
        SYNOPSYS_UNCONNECTED__230, SYNOPSYS_UNCONNECTED__231, 
        SYNOPSYS_UNCONNECTED__232, SYNOPSYS_UNCONNECTED__233, 
        SYNOPSYS_UNCONNECTED__234, SYNOPSYS_UNCONNECTED__235, 
        SYNOPSYS_UNCONNECTED__236, SYNOPSYS_UNCONNECTED__237, 
        SYNOPSYS_UNCONNECTED__238, SYNOPSYS_UNCONNECTED__239, 
        SYNOPSYS_UNCONNECTED__240, SYNOPSYS_UNCONNECTED__241, 
        SYNOPSYS_UNCONNECTED__242, SYNOPSYS_UNCONNECTED__243, 
        SYNOPSYS_UNCONNECTED__244, SYNOPSYS_UNCONNECTED__245, 
        SYNOPSYS_UNCONNECTED__246, SYNOPSYS_UNCONNECTED__247, 
        SYNOPSYS_UNCONNECTED__248, SYNOPSYS_UNCONNECTED__249, 
        SYNOPSYS_UNCONNECTED__250, SYNOPSYS_UNCONNECTED__251, 
        SYNOPSYS_UNCONNECTED__252, SYNOPSYS_UNCONNECTED__253, 
        SYNOPSYS_UNCONNECTED__254, SYNOPSYS_UNCONNECTED__255, 
        SYNOPSYS_UNCONNECTED__256, SYNOPSYS_UNCONNECTED__257, 
        SYNOPSYS_UNCONNECTED__258, SYNOPSYS_UNCONNECTED__259, 
        SYNOPSYS_UNCONNECTED__260, SYNOPSYS_UNCONNECTED__261, 
        SYNOPSYS_UNCONNECTED__262, SYNOPSYS_UNCONNECTED__263, 
        SYNOPSYS_UNCONNECTED__264, SYNOPSYS_UNCONNECTED__265, 
        SYNOPSYS_UNCONNECTED__266, SYNOPSYS_UNCONNECTED__267, 
        SYNOPSYS_UNCONNECTED__268, SYNOPSYS_UNCONNECTED__269, 
        SYNOPSYS_UNCONNECTED__270, SYNOPSYS_UNCONNECTED__271, 
        SYNOPSYS_UNCONNECTED__272, SYNOPSYS_UNCONNECTED__273, 
        SYNOPSYS_UNCONNECTED__274, SYNOPSYS_UNCONNECTED__275, 
        SYNOPSYS_UNCONNECTED__276, SYNOPSYS_UNCONNECTED__277, 
        SYNOPSYS_UNCONNECTED__278, SYNOPSYS_UNCONNECTED__279, 
        SYNOPSYS_UNCONNECTED__280, SYNOPSYS_UNCONNECTED__281, 
        SYNOPSYS_UNCONNECTED__282, SYNOPSYS_UNCONNECTED__283, 
        SYNOPSYS_UNCONNECTED__284, SYNOPSYS_UNCONNECTED__285, 
        SYNOPSYS_UNCONNECTED__286, SYNOPSYS_UNCONNECTED__287, 
        SYNOPSYS_UNCONNECTED__288, SYNOPSYS_UNCONNECTED__289, 
        SYNOPSYS_UNCONNECTED__290, SYNOPSYS_UNCONNECTED__291, 
        SYNOPSYS_UNCONNECTED__292, SYNOPSYS_UNCONNECTED__293, 
        SYNOPSYS_UNCONNECTED__294, SYNOPSYS_UNCONNECTED__295, 
        SYNOPSYS_UNCONNECTED__296, SYNOPSYS_UNCONNECTED__297, 
        SYNOPSYS_UNCONNECTED__298, SYNOPSYS_UNCONNECTED__299, 
        SYNOPSYS_UNCONNECTED__300, SYNOPSYS_UNCONNECTED__301, 
        SYNOPSYS_UNCONNECTED__302, SYNOPSYS_UNCONNECTED__303, 
        SYNOPSYS_UNCONNECTED__304, SYNOPSYS_UNCONNECTED__305, 
        SYNOPSYS_UNCONNECTED__306, SYNOPSYS_UNCONNECTED__307, 
        SYNOPSYS_UNCONNECTED__308, SYNOPSYS_UNCONNECTED__309, 
        SYNOPSYS_UNCONNECTED__310, SYNOPSYS_UNCONNECTED__311, 
        SYNOPSYS_UNCONNECTED__312, SYNOPSYS_UNCONNECTED__313, 
        SYNOPSYS_UNCONNECTED__314, SYNOPSYS_UNCONNECTED__315, 
        SYNOPSYS_UNCONNECTED__316, SYNOPSYS_UNCONNECTED__317, 
        SYNOPSYS_UNCONNECTED__318, SYNOPSYS_UNCONNECTED__319, 
        SYNOPSYS_UNCONNECTED__320, SYNOPSYS_UNCONNECTED__321, 
        SYNOPSYS_UNCONNECTED__322, SYNOPSYS_UNCONNECTED__323, 
        SYNOPSYS_UNCONNECTED__324, SYNOPSYS_UNCONNECTED__325, 
        SYNOPSYS_UNCONNECTED__326, SYNOPSYS_UNCONNECTED__327, 
        SYNOPSYS_UNCONNECTED__328, SYNOPSYS_UNCONNECTED__329, 
        SYNOPSYS_UNCONNECTED__330, SYNOPSYS_UNCONNECTED__331, 
        SYNOPSYS_UNCONNECTED__332, SYNOPSYS_UNCONNECTED__333, 
        SYNOPSYS_UNCONNECTED__334, SYNOPSYS_UNCONNECTED__335, 
        SYNOPSYS_UNCONNECTED__336, SYNOPSYS_UNCONNECTED__337, 
        SYNOPSYS_UNCONNECTED__338, SYNOPSYS_UNCONNECTED__339, 
        SYNOPSYS_UNCONNECTED__340, SYNOPSYS_UNCONNECTED__341, 
        SYNOPSYS_UNCONNECTED__342, SYNOPSYS_UNCONNECTED__343, 
        SYNOPSYS_UNCONNECTED__344, SYNOPSYS_UNCONNECTED__345, 
        SYNOPSYS_UNCONNECTED__346, SYNOPSYS_UNCONNECTED__347, 
        SYNOPSYS_UNCONNECTED__348, SYNOPSYS_UNCONNECTED__349, 
        SYNOPSYS_UNCONNECTED__350, SYNOPSYS_UNCONNECTED__351, 
        SYNOPSYS_UNCONNECTED__352, SYNOPSYS_UNCONNECTED__353, 
        SYNOPSYS_UNCONNECTED__354;

  CFD2QX2 \f01_reg[0]  ( .D(n794), .CP(clk), .CD(n919), .Q(f01[0]) );
  CFD2QX2 \f02_reg[27]  ( .D(n792), .CP(clk), .CD(n901), .Q(f02[27]) );
  CFD2QX2 \f02_reg[15]  ( .D(n784), .CP(clk), .CD(n898), .Q(f02[15]) );
  CFD2QX2 \f02_reg[11]  ( .D(n776), .CP(clk), .CD(n897), .Q(f02[11]) );
  CFD2QX2 \f02_reg[7]  ( .D(n772), .CP(clk), .CD(n896), .Q(f02[7]) );
  CFD2QX2 \f02_reg[5]  ( .D(n770), .CP(clk), .CD(n896), .Q(f02[5]) );
  CFD2QX2 \f02_reg[3]  ( .D(n766), .CP(clk), .CD(n896), .Q(f02[3]) );
  CFD2QX2 \f03_reg[18]  ( .D(n750), .CP(clk), .CD(n888), .Q(f03[18]) );
  CFD2QX2 \f03_reg[17]  ( .D(n748), .CP(clk), .CD(n888), .Q(f03[17]) );
  CFD2QX2 \f03_reg[14]  ( .D(n746), .CP(clk), .CD(n887), .Q(f03[14]) );
  CFD2QX2 \f03_reg[12]  ( .D(n744), .CP(clk), .CD(n887), .Q(f03[12]) );
  CFD2QX2 \f03_reg[10]  ( .D(n742), .CP(clk), .CD(n886), .Q(f03[10]) );
  CFD2QX2 \f03_reg[6]  ( .D(n740), .CP(clk), .CD(n886), .Q(f03[6]) );
  CFD2QX2 \f03_reg[0]  ( .D(n732), .CP(clk), .CD(n885), .Q(f03[0]) );
  CFD2QX2 \f11_reg[20]  ( .D(n728), .CP(clk), .CD(n916), .Q(f11[20]) );
  CFD2QX2 \f11_reg[2]  ( .D(n724), .CP(clk), .CD(n915), .Q(f11[2]) );
  CFD2QX2 \f12_reg[29]  ( .D(s12[29]), .CP(clk), .CD(n919), .Q(f12[29]) );
  CFD2QX2 \f12_reg[18]  ( .D(s12[18]), .CP(clk), .CD(n918), .Q(f12[18]) );
  CFD2QX2 \f12_reg[14]  ( .D(s12[14]), .CP(clk), .CD(n918), .Q(f12[14]) );
  CFD2QX2 \f12_reg[12]  ( .D(s12[12]), .CP(clk), .CD(n918), .Q(f12[12]) );
  CFD2QX2 \f12_reg[10]  ( .D(s12[10]), .CP(clk), .CD(n918), .Q(f12[10]) );
  CFD2QX2 \f12_reg[4]  ( .D(s12[4]), .CP(clk), .CD(n917), .Q(f12[4]) );
  CFD2QX2 \f12_reg[3]  ( .D(s12[3]), .CP(clk), .CD(n917), .Q(f12[3]) );
  CFD2QX2 \f13_reg[27]  ( .D(n722), .CP(clk), .CD(n901), .Q(f13[27]) );
  CFD2QX2 \f13_reg[25]  ( .D(n719), .CP(clk), .CD(n901), .Q(f13[25]) );
  CFD2QX2 \f13_reg[18]  ( .D(n708), .CP(clk), .CD(n899), .Q(f13[18]) );
  CFD2QX2 \f13_reg[16]  ( .D(n706), .CP(clk), .CD(n898), .Q(f13[16]) );
  CFD2QX2 \f13_reg[14]  ( .D(n705), .CP(clk), .CD(n898), .Q(f13[14]) );
  CFD2QX2 \f13_reg[12]  ( .D(n703), .CP(clk), .CD(n898), .Q(f13[12]) );
  calc_DW01_add_6 add_208 ( .A(f16), .B(f17), .CI(1'b0), .SUM(s27) );
  calc_DW01_add_7 add_232 ( .A(f51), .B(f52), .CI(1'b0), .SUM(res_temp) );
  calc_DW01_add_8 add_227 ( .A(f41), .B(f42), .CI(1'b0), .SUM(s51) );
  calc_DW01_add_9 add_223 ( .A(f33), .B({f34[31:2], 1'b0, f34[0]}), .CI(1'b0), 
        .SUM(s43) );
  calc_DW01_add_10 add_215 ( .A(f24), .B(f22), .CI(1'b0), .SUM(s33) );
  calc_DW01_add_11 add_214 ( .A(f26), .B(f27), .CI(1'b0), .SUM(s32) );
  calc_DW_mult_uns_11 mult_205 ( .a({f12[31:20], n828, f12[18:3], n123, 1'b0, 
        f12[0]}), .b(f17), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, s24}) );
  calc_DW_mult_uns_12 mult_204 ( .a({f12[31:3], n123, 1'b0, f12[0]}), .b({
        f11[31:22], n835, f11[20], n829, f11[18:4], n128, f11[2:0]}), 
        .product({SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, s23}) );
  calc_DW_mult_uns_13 mult_203 ( .a(f11), .b({f13[31:20], n832, f13[18], n125, 
        f13[16:6], n837, f13[4], n839, f13[2:0]}), .product({
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, s22}) );
  calc_DW_mult_uns_14 mult_207 ( .a(f13), .b({f14[31:2], 1'b0, f14[0]}), 
        .product({SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, s26}) );
  calc_DW_mult_uns_15 mult_198 ( .a(f02), .b(f03), .product({
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, s17}) );
  calc_DW_mult_uns_16 mult_197 ( .a(f01), .b(f03), .product({
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, 
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        SYNOPSYS_UNCONNECTED__174, SYNOPSYS_UNCONNECTED__175, 
        SYNOPSYS_UNCONNECTED__176, SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, 
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        SYNOPSYS_UNCONNECTED__184, SYNOPSYS_UNCONNECTED__185, 
        SYNOPSYS_UNCONNECTED__186, SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, s16}) );
  calc_DW_mult_uns_17 mult_213 ( .a(f23), .b(f21), .product({
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, 
        SYNOPSYS_UNCONNECTED__202, SYNOPSYS_UNCONNECTED__203, 
        SYNOPSYS_UNCONNECTED__204, SYNOPSYS_UNCONNECTED__205, 
        SYNOPSYS_UNCONNECTED__206, SYNOPSYS_UNCONNECTED__207, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, 
        SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213, 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        SYNOPSYS_UNCONNECTED__216, SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, 
        SYNOPSYS_UNCONNECTED__222, SYNOPSYS_UNCONNECTED__223, s31}) );
  calc_DW_mult_uns_18 mult_221 ( .a({f31[31:13], n830, f31[11:0]}), .b(f30), 
        .product({SYNOPSYS_UNCONNECTED__224, SYNOPSYS_UNCONNECTED__225, 
        SYNOPSYS_UNCONNECTED__226, SYNOPSYS_UNCONNECTED__227, 
        SYNOPSYS_UNCONNECTED__228, SYNOPSYS_UNCONNECTED__229, 
        SYNOPSYS_UNCONNECTED__230, SYNOPSYS_UNCONNECTED__231, 
        SYNOPSYS_UNCONNECTED__232, SYNOPSYS_UNCONNECTED__233, 
        SYNOPSYS_UNCONNECTED__234, SYNOPSYS_UNCONNECTED__235, 
        SYNOPSYS_UNCONNECTED__236, SYNOPSYS_UNCONNECTED__237, 
        SYNOPSYS_UNCONNECTED__238, SYNOPSYS_UNCONNECTED__239, 
        SYNOPSYS_UNCONNECTED__240, SYNOPSYS_UNCONNECTED__241, 
        SYNOPSYS_UNCONNECTED__242, SYNOPSYS_UNCONNECTED__243, 
        SYNOPSYS_UNCONNECTED__244, SYNOPSYS_UNCONNECTED__245, 
        SYNOPSYS_UNCONNECTED__246, SYNOPSYS_UNCONNECTED__247, 
        SYNOPSYS_UNCONNECTED__248, SYNOPSYS_UNCONNECTED__249, 
        SYNOPSYS_UNCONNECTED__250, SYNOPSYS_UNCONNECTED__251, 
        SYNOPSYS_UNCONNECTED__252, SYNOPSYS_UNCONNECTED__253, 
        SYNOPSYS_UNCONNECTED__254, SYNOPSYS_UNCONNECTED__255, s41}) );
  calc_DW_mult_uns_19 mult_196 ( .a(f03), .b({f03[31:1], n264}), .product({
        SYNOPSYS_UNCONNECTED__256, SYNOPSYS_UNCONNECTED__257, 
        SYNOPSYS_UNCONNECTED__258, SYNOPSYS_UNCONNECTED__259, 
        SYNOPSYS_UNCONNECTED__260, SYNOPSYS_UNCONNECTED__261, 
        SYNOPSYS_UNCONNECTED__262, SYNOPSYS_UNCONNECTED__263, 
        SYNOPSYS_UNCONNECTED__264, SYNOPSYS_UNCONNECTED__265, 
        SYNOPSYS_UNCONNECTED__266, SYNOPSYS_UNCONNECTED__267, 
        SYNOPSYS_UNCONNECTED__268, SYNOPSYS_UNCONNECTED__269, 
        SYNOPSYS_UNCONNECTED__270, SYNOPSYS_UNCONNECTED__271, 
        SYNOPSYS_UNCONNECTED__272, SYNOPSYS_UNCONNECTED__273, 
        SYNOPSYS_UNCONNECTED__274, SYNOPSYS_UNCONNECTED__275, 
        SYNOPSYS_UNCONNECTED__276, SYNOPSYS_UNCONNECTED__277, 
        SYNOPSYS_UNCONNECTED__278, SYNOPSYS_UNCONNECTED__279, 
        SYNOPSYS_UNCONNECTED__280, SYNOPSYS_UNCONNECTED__281, 
        SYNOPSYS_UNCONNECTED__282, SYNOPSYS_UNCONNECTED__283, 
        SYNOPSYS_UNCONNECTED__284, SYNOPSYS_UNCONNECTED__285, 
        SYNOPSYS_UNCONNECTED__286, SYNOPSYS_UNCONNECTED__287, s15[31:2], 
        SYNOPSYS_UNCONNECTED__288, s15[0]}) );
  calc_DW_mult_uns_20 mult_195 ( .a({f02[31:16], n124, f02[14:0]}), .b({
        f02[31:16], n124, f02[14:1], n693}), .product({
        SYNOPSYS_UNCONNECTED__289, SYNOPSYS_UNCONNECTED__290, 
        SYNOPSYS_UNCONNECTED__291, SYNOPSYS_UNCONNECTED__292, 
        SYNOPSYS_UNCONNECTED__293, SYNOPSYS_UNCONNECTED__294, 
        SYNOPSYS_UNCONNECTED__295, SYNOPSYS_UNCONNECTED__296, 
        SYNOPSYS_UNCONNECTED__297, SYNOPSYS_UNCONNECTED__298, 
        SYNOPSYS_UNCONNECTED__299, SYNOPSYS_UNCONNECTED__300, 
        SYNOPSYS_UNCONNECTED__301, SYNOPSYS_UNCONNECTED__302, 
        SYNOPSYS_UNCONNECTED__303, SYNOPSYS_UNCONNECTED__304, 
        SYNOPSYS_UNCONNECTED__305, SYNOPSYS_UNCONNECTED__306, 
        SYNOPSYS_UNCONNECTED__307, SYNOPSYS_UNCONNECTED__308, 
        SYNOPSYS_UNCONNECTED__309, SYNOPSYS_UNCONNECTED__310, 
        SYNOPSYS_UNCONNECTED__311, SYNOPSYS_UNCONNECTED__312, 
        SYNOPSYS_UNCONNECTED__313, SYNOPSYS_UNCONNECTED__314, 
        SYNOPSYS_UNCONNECTED__315, SYNOPSYS_UNCONNECTED__316, 
        SYNOPSYS_UNCONNECTED__317, SYNOPSYS_UNCONNECTED__318, 
        SYNOPSYS_UNCONNECTED__319, SYNOPSYS_UNCONNECTED__320, s14[31:2], 
        SYNOPSYS_UNCONNECTED__321, s14[0]}) );
  calc_DW_mult_uns_21 mult_193 ( .a({f01[31:16], n833, f01[14], n127, 
        f01[12:6], n126, f01[4:0]}), .b({f01[31:14], n127, f01[12:6], n126, 
        f01[4:1], n121}), .product({SYNOPSYS_UNCONNECTED__322, 
        SYNOPSYS_UNCONNECTED__323, SYNOPSYS_UNCONNECTED__324, 
        SYNOPSYS_UNCONNECTED__325, SYNOPSYS_UNCONNECTED__326, 
        SYNOPSYS_UNCONNECTED__327, SYNOPSYS_UNCONNECTED__328, 
        SYNOPSYS_UNCONNECTED__329, SYNOPSYS_UNCONNECTED__330, 
        SYNOPSYS_UNCONNECTED__331, SYNOPSYS_UNCONNECTED__332, 
        SYNOPSYS_UNCONNECTED__333, SYNOPSYS_UNCONNECTED__334, 
        SYNOPSYS_UNCONNECTED__335, SYNOPSYS_UNCONNECTED__336, 
        SYNOPSYS_UNCONNECTED__337, SYNOPSYS_UNCONNECTED__338, 
        SYNOPSYS_UNCONNECTED__339, SYNOPSYS_UNCONNECTED__340, 
        SYNOPSYS_UNCONNECTED__341, SYNOPSYS_UNCONNECTED__342, 
        SYNOPSYS_UNCONNECTED__343, SYNOPSYS_UNCONNECTED__344, 
        SYNOPSYS_UNCONNECTED__345, SYNOPSYS_UNCONNECTED__346, 
        SYNOPSYS_UNCONNECTED__347, SYNOPSYS_UNCONNECTED__348, 
        SYNOPSYS_UNCONNECTED__349, SYNOPSYS_UNCONNECTED__350, 
        SYNOPSYS_UNCONNECTED__351, SYNOPSYS_UNCONNECTED__352, 
        SYNOPSYS_UNCONNECTED__353, s12[31:2], SYNOPSYS_UNCONNECTED__354, 
        s12[0]}) );
  CFD2QX1 \f13_reg[5]  ( .D(n600), .CP(clk), .CD(n896), .Q(f13[5]) );
  CFD2QXL \f15_reg[27]  ( .D(s15[27]), .CP(clk), .CD(n862), .Q(f15[27]) );
  CFD2QXL \f21_reg[15]  ( .D(f11[15]), .CP(clk), .CD(n911), .Q(f21[15]) );
  CFD2QX1 \f12_reg[19]  ( .D(s12[19]), .CP(clk), .CD(n918), .Q(f12[19]) );
  CFD2QXL \f21_reg[3]  ( .D(n596), .CP(clk), .CD(n910), .Q(f21[3]) );
  CFD2QX1 \f13_reg[15]  ( .D(n124), .CP(clk), .CD(n898), .Q(f13[15]) );
  CFD2QX1 \f12_reg[21]  ( .D(s12[21]), .CP(clk), .CD(n919), .Q(f12[21]) );
  CFD2QX1 \f11_reg[13]  ( .D(n593), .CP(clk), .CD(n915), .Q(f11[13]) );
  CFD2QX1 \f13_reg[13]  ( .D(n591), .CP(clk), .CD(n898), .Q(f13[13]) );
  CFD2QX4 \f11_reg[12]  ( .D(n588), .CP(clk), .CD(n915), .Q(f11[12]) );
  CFD2QX1 \f11_reg[11]  ( .D(n589), .CP(clk), .CD(n915), .Q(f11[11]) );
  CFD2QX1 \f13_reg[11]  ( .D(n586), .CP(clk), .CD(n897), .Q(f13[11]) );
  CFD2QX1 \f23_reg[5]  ( .D(s23[5]), .CP(clk), .CD(n912), .Q(f23[5]) );
  CFD2QX1 \f13_reg[3]  ( .D(n584), .CP(clk), .CD(n895), .Q(f13[3]) );
  CFD2QX1 \f13_reg[7]  ( .D(n582), .CP(clk), .CD(n896), .Q(f13[7]) );
  CFD2QX1 \f23_reg[13]  ( .D(s23[13]), .CP(clk), .CD(n913), .Q(f23[13]) );
  CFD2QX1 \f01_reg[13]  ( .D(n579), .CP(clk), .CD(n921), .Q(f01[13]) );
  CFD2QX1 \f21_reg[19]  ( .D(n829), .CP(clk), .CD(n911), .Q(f21[19]) );
  CFD2QX1 \f31_reg[7]  ( .D(s31[7]), .CP(clk), .CD(n908), .Q(f31[7]) );
  CFD2QX1 \f31_reg[5]  ( .D(s31[5]), .CP(clk), .CD(n907), .Q(f31[5]) );
  CFD2QX1 \f13_reg[1]  ( .D(n575), .CP(clk), .CD(n895), .Q(f13[1]) );
  CFD2QXL \f31_reg[31]  ( .D(s31[31]), .CP(clk), .CD(n909), .Q(f31[31]) );
  CFD2QX1 \f31_reg[9]  ( .D(s31[9]), .CP(clk), .CD(n908), .Q(f31[9]) );
  CFD2QX1 \f01_reg[19]  ( .D(n573), .CP(clk), .CD(n922), .Q(f01[19]) );
  CFD2QX4 \f12_reg[27]  ( .D(s12[27]), .CP(clk), .CD(n919), .Q(f12[27]) );
  CFD2QX1 \f23_reg[15]  ( .D(s23[15]), .CP(clk), .CD(n913), .Q(f23[15]) );
  CFD2QX1 \f02_reg[21]  ( .D(n571), .CP(clk), .CD(n900), .Q(f02[21]) );
  CFD2QX1 \f13_reg[17]  ( .D(n568), .CP(clk), .CD(n899), .Q(f13[17]) );
  CFD2QX1 \f23_reg[9]  ( .D(s23[9]), .CP(clk), .CD(n913), .Q(f23[9]) );
  CFD2QX1 \f21_reg[17]  ( .D(n566), .CP(clk), .CD(n911), .Q(f21[17]) );
  CFD2QXL \captA_reg[19]  ( .D(n105), .CP(clk), .CD(n922), .Q(captA[19]) );
  CFD2QXL \captA_reg[13]  ( .D(n99), .CP(clk), .CD(n921), .Q(captA[13]) );
  CFD2QXL \captB_reg[21]  ( .D(n75), .CP(clk), .CD(n900), .Q(captB[21]) );
  CFD2QXL \captB_reg[6]  ( .D(n60), .CP(clk), .CD(n896), .Q(captB[6]) );
  CFD2QXL \captC_reg[16]  ( .D(n38), .CP(clk), .CD(n887), .Q(captC[16]) );
  CFD2QXL \captC_reg[15]  ( .D(n37), .CP(clk), .CD(n887), .Q(captC[15]) );
  CFD2QXL \captC_reg[9]  ( .D(n31), .CP(clk), .CD(n886), .Q(captC[9]) );
  CFD2QXL \captC_reg[8]  ( .D(n30), .CP(clk), .CD(n886), .Q(captC[8]) );
  CFD2QXL \captC_reg[5]  ( .D(n27), .CP(clk), .CD(n886), .Q(captC[5]) );
  CFD2QXL \captA_reg[31]  ( .D(n117), .CP(clk), .CD(n924), .Q(captA[31]) );
  CFD2QXL \captA_reg[30]  ( .D(n116), .CP(clk), .CD(n924), .Q(captA[30]) );
  CFD2QXL \captA_reg[29]  ( .D(n115), .CP(clk), .CD(n924), .Q(captA[29]) );
  CFD2QXL \captA_reg[28]  ( .D(n114), .CP(clk), .CD(n924), .Q(captA[28]) );
  CFD2QXL \captA_reg[27]  ( .D(n113), .CP(clk), .CD(n924), .Q(captA[27]) );
  CFD2QXL \captA_reg[26]  ( .D(n112), .CP(clk), .CD(n923), .Q(captA[26]) );
  CFD2QXL \captA_reg[25]  ( .D(n111), .CP(clk), .CD(n923), .Q(captA[25]) );
  CFD2QXL \captA_reg[24]  ( .D(n110), .CP(clk), .CD(n923), .Q(captA[24]) );
  CFD2QXL \captA_reg[23]  ( .D(n109), .CP(clk), .CD(n923), .Q(captA[23]) );
  CFD2QXL \captA_reg[22]  ( .D(n108), .CP(clk), .CD(n923), .Q(captA[22]) );
  CFD2QXL \captA_reg[21]  ( .D(n107), .CP(clk), .CD(n923), .Q(captA[21]) );
  CFD2QXL \captA_reg[20]  ( .D(n106), .CP(clk), .CD(n923), .Q(captA[20]) );
  CFD2QXL \captA_reg[18]  ( .D(n104), .CP(clk), .CD(n922), .Q(captA[18]) );
  CFD2QXL \captA_reg[17]  ( .D(n103), .CP(clk), .CD(n922), .Q(captA[17]) );
  CFD2QXL \captA_reg[16]  ( .D(n102), .CP(clk), .CD(n922), .Q(captA[16]) );
  CFD2QXL \captA_reg[15]  ( .D(n101), .CP(clk), .CD(n922), .Q(captA[15]) );
  CFD2QXL \captA_reg[14]  ( .D(n100), .CP(clk), .CD(n922), .Q(captA[14]) );
  CFD2QXL \captA_reg[12]  ( .D(n98), .CP(clk), .CD(n921), .Q(captA[12]) );
  CFD2QXL \captA_reg[11]  ( .D(n97), .CP(clk), .CD(n921), .Q(captA[11]) );
  CFD2QXL \captA_reg[10]  ( .D(n96), .CP(clk), .CD(n921), .Q(captA[10]) );
  CFD2QXL \captA_reg[9]  ( .D(n95), .CP(clk), .CD(n921), .Q(captA[9]) );
  CFD2QXL \captA_reg[8]  ( .D(n94), .CP(clk), .CD(n921), .Q(captA[8]) );
  CFD2QXL \captA_reg[7]  ( .D(n93), .CP(clk), .CD(n921), .Q(captA[7]) );
  CFD2QXL \captA_reg[6]  ( .D(n92), .CP(clk), .CD(n920), .Q(captA[6]) );
  CFD2QXL \captA_reg[5]  ( .D(n91), .CP(clk), .CD(n920), .Q(captA[5]) );
  CFD2QXL \captA_reg[4]  ( .D(n90), .CP(clk), .CD(n920), .Q(captA[4]) );
  CFD2QXL \captA_reg[3]  ( .D(n89), .CP(clk), .CD(n920), .Q(captA[3]) );
  CFD2QXL \captA_reg[2]  ( .D(n88), .CP(clk), .CD(n920), .Q(captA[2]) );
  CFD2QXL \captA_reg[1]  ( .D(n87), .CP(clk), .CD(n920), .Q(captA[1]) );
  CFD2QXL \captA_reg[0]  ( .D(n86), .CP(clk), .CD(n919), .Q(captA[0]) );
  CFD2QXL \captB_reg[31]  ( .D(n85), .CP(clk), .CD(n902), .Q(captB[31]) );
  CFD2QXL \captB_reg[30]  ( .D(n84), .CP(clk), .CD(n902), .Q(captB[30]) );
  CFD2QXL \captB_reg[29]  ( .D(n83), .CP(clk), .CD(n902), .Q(captB[29]) );
  CFD2QXL \captB_reg[28]  ( .D(n82), .CP(clk), .CD(n901), .Q(captB[28]) );
  CFD2QXL \captB_reg[27]  ( .D(n81), .CP(clk), .CD(n901), .Q(captB[27]) );
  CFD2QXL \captB_reg[26]  ( .D(n80), .CP(clk), .CD(n901), .Q(captB[26]) );
  CFD2QXL \captB_reg[25]  ( .D(n79), .CP(clk), .CD(n901), .Q(captB[25]) );
  CFD2QXL \captB_reg[24]  ( .D(n78), .CP(clk), .CD(n900), .Q(captB[24]) );
  CFD2QXL \captB_reg[23]  ( .D(n77), .CP(clk), .CD(n900), .Q(captB[23]) );
  CFD2QXL \captB_reg[22]  ( .D(n76), .CP(clk), .CD(n900), .Q(captB[22]) );
  CFD2QXL \captB_reg[20]  ( .D(n74), .CP(clk), .CD(n900), .Q(captB[20]) );
  CFD2QXL \captB_reg[19]  ( .D(n73), .CP(clk), .CD(n899), .Q(captB[19]) );
  CFD2QXL \captB_reg[18]  ( .D(n72), .CP(clk), .CD(n899), .Q(captB[18]) );
  CFD2QXL \captB_reg[17]  ( .D(n71), .CP(clk), .CD(n899), .Q(captB[17]) );
  CFD2QXL \captB_reg[16]  ( .D(n70), .CP(clk), .CD(n899), .Q(captB[16]) );
  CFD2QXL \captB_reg[15]  ( .D(n69), .CP(clk), .CD(n898), .Q(captB[15]) );
  CFD2QXL \captB_reg[14]  ( .D(n68), .CP(clk), .CD(n898), .Q(captB[14]) );
  CFD2QXL \captB_reg[13]  ( .D(n67), .CP(clk), .CD(n898), .Q(captB[13]) );
  CFD2QXL \captB_reg[12]  ( .D(n66), .CP(clk), .CD(n898), .Q(captB[12]) );
  CFD2QXL \captB_reg[11]  ( .D(n65), .CP(clk), .CD(n897), .Q(captB[11]) );
  CFD2QXL \captB_reg[10]  ( .D(n64), .CP(clk), .CD(n897), .Q(captB[10]) );
  CFD2QXL \captB_reg[9]  ( .D(n63), .CP(clk), .CD(n897), .Q(captB[9]) );
  CFD2QXL \captB_reg[8]  ( .D(n62), .CP(clk), .CD(n897), .Q(captB[8]) );
  CFD2QXL \captB_reg[7]  ( .D(n61), .CP(clk), .CD(n897), .Q(captB[7]) );
  CFD2QXL \captB_reg[5]  ( .D(n59), .CP(clk), .CD(n896), .Q(captB[5]) );
  CFD2QXL \captB_reg[4]  ( .D(n58), .CP(clk), .CD(n896), .Q(captB[4]) );
  CFD2QXL \captB_reg[3]  ( .D(n57), .CP(clk), .CD(n896), .Q(captB[3]) );
  CFD2QXL \captB_reg[2]  ( .D(n56), .CP(clk), .CD(n895), .Q(captB[2]) );
  CFD2QXL \captB_reg[1]  ( .D(n55), .CP(clk), .CD(n895), .Q(captB[1]) );
  CFD2QXL \captB_reg[0]  ( .D(n54), .CP(clk), .CD(n895), .Q(captB[0]) );
  CFD2QXL \captC_reg[31]  ( .D(n53), .CP(clk), .CD(n890), .Q(captC[31]) );
  CFD2QXL \captC_reg[30]  ( .D(n52), .CP(clk), .CD(n890), .Q(captC[30]) );
  CFD2QXL \captC_reg[29]  ( .D(n51), .CP(clk), .CD(n889), .Q(captC[29]) );
  CFD2QXL \captC_reg[28]  ( .D(n50), .CP(clk), .CD(n889), .Q(captC[28]) );
  CFD2QXL \captC_reg[27]  ( .D(n49), .CP(clk), .CD(n889), .Q(captC[27]) );
  CFD2QXL \captC_reg[26]  ( .D(n48), .CP(clk), .CD(n889), .Q(captC[26]) );
  CFD2QXL \captC_reg[25]  ( .D(n47), .CP(clk), .CD(n889), .Q(captC[25]) );
  CFD2QXL \captC_reg[24]  ( .D(n46), .CP(clk), .CD(n889), .Q(captC[24]) );
  CFD2QXL \captC_reg[23]  ( .D(n45), .CP(clk), .CD(n889), .Q(captC[23]) );
  CFD2QXL \captC_reg[22]  ( .D(n44), .CP(clk), .CD(n888), .Q(captC[22]) );
  CFD2QXL \captC_reg[21]  ( .D(n43), .CP(clk), .CD(n888), .Q(captC[21]) );
  CFD2QXL \captC_reg[20]  ( .D(n42), .CP(clk), .CD(n888), .Q(captC[20]) );
  CFD2QXL \captC_reg[19]  ( .D(n41), .CP(clk), .CD(n888), .Q(captC[19]) );
  CFD2QXL \captC_reg[18]  ( .D(n40), .CP(clk), .CD(n888), .Q(captC[18]) );
  CFD2QXL \captC_reg[17]  ( .D(n39), .CP(clk), .CD(n888), .Q(captC[17]) );
  CFD2QXL \captC_reg[14]  ( .D(n36), .CP(clk), .CD(n887), .Q(captC[14]) );
  CFD2QXL \captC_reg[13]  ( .D(n35), .CP(clk), .CD(n887), .Q(captC[13]) );
  CFD2QXL \captC_reg[12]  ( .D(n34), .CP(clk), .CD(n887), .Q(captC[12]) );
  CFD2QXL \captC_reg[11]  ( .D(n33), .CP(clk), .CD(n887), .Q(captC[11]) );
  CFD2QXL \captC_reg[10]  ( .D(n32), .CP(clk), .CD(n887), .Q(captC[10]) );
  CFD2QXL \captC_reg[7]  ( .D(n29), .CP(clk), .CD(n886), .Q(captC[7]) );
  CFD2QXL \captC_reg[6]  ( .D(n28), .CP(clk), .CD(n886), .Q(captC[6]) );
  CFD2QXL \captC_reg[4]  ( .D(n26), .CP(clk), .CD(n886), .Q(captC[4]) );
  CFD2QXL \captC_reg[3]  ( .D(n25), .CP(clk), .CD(n885), .Q(captC[3]) );
  CFD2QXL \captC_reg[2]  ( .D(n24), .CP(clk), .CD(n885), .Q(captC[2]) );
  CFD2QXL \captC_reg[1]  ( .D(n23), .CP(clk), .CD(n885), .Q(captC[1]) );
  CFD2QXL \captC_reg[0]  ( .D(n22), .CP(clk), .CD(n885), .Q(captC[0]) );
  CFD2QXL \f24_reg[30]  ( .D(s24[30]), .CP(clk), .CD(n870), .Q(f24[30]) );
  CFD2QXL \f24_reg[29]  ( .D(s24[29]), .CP(clk), .CD(n870), .Q(f24[29]) );
  CFD2QXL \f24_reg[28]  ( .D(s24[28]), .CP(clk), .CD(n870), .Q(f24[28]) );
  CFD2QXL \f26_reg[30]  ( .D(s26[30]), .CP(clk), .CD(n892), .Q(f26[30]) );
  CFD2QXL \f26_reg[29]  ( .D(s26[29]), .CP(clk), .CD(n892), .Q(f26[29]) );
  CFD2QXL \f26_reg[28]  ( .D(s26[28]), .CP(clk), .CD(n892), .Q(f26[28]) );
  CFD2QXL \f33_reg[30]  ( .D(s33[30]), .CP(clk), .CD(n865), .Q(f33[30]) );
  CFD2QXL \f33_reg[29]  ( .D(s33[29]), .CP(clk), .CD(n865), .Q(f33[29]) );
  CFD2QXL \f33_reg[28]  ( .D(s33[28]), .CP(clk), .CD(n865), .Q(f33[28]) );
  CFD2QXL \f41_reg[30]  ( .D(s41[30]), .CP(clk), .CD(n904), .Q(f41[30]) );
  CFD2QXL \f41_reg[29]  ( .D(s41[29]), .CP(clk), .CD(n904), .Q(f41[29]) );
  CFD2QXL \f41_reg[28]  ( .D(s41[28]), .CP(clk), .CD(n904), .Q(f41[28]) );
  CFD2QXL \f51_reg[28]  ( .D(s51[28]), .CP(clk), .CD(n872), .Q(f51[28]) );
  CFD2QXL \f51_reg[29]  ( .D(s51[29]), .CP(clk), .CD(n872), .Q(f51[29]) );
  CFD2QXL \f51_reg[30]  ( .D(s51[30]), .CP(clk), .CD(n872), .Q(f51[30]) );
  CFD2QXL \f16_reg[30]  ( .D(s16[30]), .CP(clk), .CD(n885), .Q(f16[30]) );
  CFD2QXL \f16_reg[29]  ( .D(s16[29]), .CP(clk), .CD(n885), .Q(f16[29]) );
  CFD2QXL \f16_reg[28]  ( .D(s16[28]), .CP(clk), .CD(n885), .Q(f16[28]) );
  CFD2QXL \f16_reg[27]  ( .D(s16[27]), .CP(clk), .CD(n885), .Q(f16[27]) );
  CFD2QXL \f22_reg[30]  ( .D(s22[30]), .CP(clk), .CD(n868), .Q(f22[30]) );
  CFD2QXL \f22_reg[29]  ( .D(s22[29]), .CP(clk), .CD(n867), .Q(f22[29]) );
  CFD2QXL \f22_reg[28]  ( .D(s22[28]), .CP(clk), .CD(n867), .Q(f22[28]) );
  CFD2QXL \f27_reg[30]  ( .D(s27[30]), .CP(clk), .CD(n880), .Q(f27[30]) );
  CFD2QXL \f27_reg[29]  ( .D(s27[29]), .CP(clk), .CD(n880), .Q(f27[29]) );
  CFD2QXL \f27_reg[28]  ( .D(s27[28]), .CP(clk), .CD(n880), .Q(f27[28]) );
  CFD2QXL \f34_reg[30]  ( .D(n551), .CP(clk), .CD(n862), .Q(f34[30]) );
  CFD2QXL \f34_reg[29]  ( .D(n549), .CP(clk), .CD(n862), .Q(f34[29]) );
  CFD2QXL \f34_reg[28]  ( .D(n547), .CP(clk), .CD(n862), .Q(f34[28]) );
  CFD2QXL \f42_reg[30]  ( .D(n545), .CP(clk), .CD(n877), .Q(f42[30]) );
  CFD2QXL \f42_reg[29]  ( .D(n543), .CP(clk), .CD(n877), .Q(f42[29]) );
  CFD2QXL \f42_reg[28]  ( .D(n541), .CP(clk), .CD(n877), .Q(f42[28]) );
  CFD2QXL \f52_reg[30]  ( .D(n539), .CP(clk), .CD(n855), .Q(f52[30]) );
  CFD2QXL \f52_reg[29]  ( .D(n537), .CP(clk), .CD(n855), .Q(f52[29]) );
  CFD2QXL \f52_reg[28]  ( .D(n535), .CP(clk), .CD(n855), .Q(f52[28]) );
  CFD2QXL \f24_reg[31]  ( .D(s24[31]), .CP(clk), .CD(n870), .Q(f24[31]) );
  CFD2QXL \f26_reg[31]  ( .D(s26[31]), .CP(clk), .CD(n892), .Q(f26[31]) );
  CFD2QXL \f33_reg[31]  ( .D(s33[31]), .CP(clk), .CD(n865), .Q(f33[31]) );
  CFD2QXL \f41_reg[31]  ( .D(s41[31]), .CP(clk), .CD(n905), .Q(f41[31]) );
  CFD2QXL \f51_reg[31]  ( .D(s51[31]), .CP(clk), .CD(n873), .Q(f51[31]) );
  CFD2QXL \f26_reg[27]  ( .D(s26[27]), .CP(clk), .CD(n892), .Q(f26[27]) );
  CFD2QXL \f41_reg[27]  ( .D(s41[27]), .CP(clk), .CD(n904), .Q(f41[27]) );
  CFD2QXL \f51_reg[27]  ( .D(s51[27]), .CP(clk), .CD(n872), .Q(f51[27]) );
  CFD2QXL \f16_reg[31]  ( .D(s16[31]), .CP(clk), .CD(n885), .Q(f16[31]) );
  CFD2QXL \f22_reg[31]  ( .D(s22[31]), .CP(clk), .CD(n868), .Q(f22[31]) );
  CFD2QXL \f27_reg[31]  ( .D(s27[31]), .CP(clk), .CD(n880), .Q(f27[31]) );
  CFD2QXL \f34_reg[31]  ( .D(n533), .CP(clk), .CD(n863), .Q(f34[31]) );
  CFD2QXL \f42_reg[31]  ( .D(n531), .CP(clk), .CD(n877), .Q(f42[31]) );
  CFD2QXL \f52_reg[31]  ( .D(n529), .CP(clk), .CD(n855), .Q(f52[31]) );
  CFD2QXL \seen_reg[1]  ( .D(seen_d[1]), .CP(clk), .CD(n925), .Q(stopB) );
  CFD2QXL \seen_reg[0]  ( .D(seen_d[0]), .CP(clk), .CD(n924), .Q(stopC) );
  CFD2QXL \seen_reg[2]  ( .D(seen_d[2]), .CP(clk), .CD(n925), .Q(stopA) );
  CFD2QXL \f30_reg[31]  ( .D(n527), .CP(clk), .CD(n907), .Q(f30[31]) );
  CFD2QXL \f03_reg[31]  ( .D(n526), .CP(clk), .CD(n890), .Q(f03[31]) );
  CFD2QXL \f14_reg[31]  ( .D(s14[31]), .CP(clk), .CD(n895), .Q(f14[31]) );
  CFD2QXL \f24_reg[27]  ( .D(s24[27]), .CP(clk), .CD(n870), .Q(f24[27]) );
  CFD2QXL \f24_reg[26]  ( .D(s24[26]), .CP(clk), .CD(n870), .Q(f24[26]) );
  CFD2QXL \f24_reg[25]  ( .D(s24[25]), .CP(clk), .CD(n870), .Q(f24[25]) );
  CFD2QXL \f24_reg[24]  ( .D(s24[24]), .CP(clk), .CD(n870), .Q(f24[24]) );
  CFD2QXL \f24_reg[23]  ( .D(s24[23]), .CP(clk), .CD(n869), .Q(f24[23]) );
  CFD2QXL \f24_reg[22]  ( .D(s24[22]), .CP(clk), .CD(n869), .Q(f24[22]) );
  CFD2QXL \f24_reg[21]  ( .D(s24[21]), .CP(clk), .CD(n869), .Q(f24[21]) );
  CFD2QXL \f24_reg[20]  ( .D(s24[20]), .CP(clk), .CD(n869), .Q(f24[20]) );
  CFD2QXL \f26_reg[26]  ( .D(s26[26]), .CP(clk), .CD(n892), .Q(f26[26]) );
  CFD2QXL \f26_reg[25]  ( .D(s26[25]), .CP(clk), .CD(n892), .Q(f26[25]) );
  CFD2QXL \f26_reg[24]  ( .D(s26[24]), .CP(clk), .CD(n892), .Q(f26[24]) );
  CFD2QXL \f26_reg[23]  ( .D(s26[23]), .CP(clk), .CD(n892), .Q(f26[23]) );
  CFD2QXL \f26_reg[22]  ( .D(s26[22]), .CP(clk), .CD(n892), .Q(f26[22]) );
  CFD2QXL \f26_reg[21]  ( .D(s26[21]), .CP(clk), .CD(n891), .Q(f26[21]) );
  CFD2QXL \f26_reg[20]  ( .D(s26[20]), .CP(clk), .CD(n891), .Q(f26[20]) );
  CFD2QXL \f26_reg[19]  ( .D(s26[19]), .CP(clk), .CD(n891), .Q(f26[19]) );
  CFD2QXL \f26_reg[18]  ( .D(s26[18]), .CP(clk), .CD(n891), .Q(f26[18]) );
  CFD2QXL \f33_reg[27]  ( .D(s33[27]), .CP(clk), .CD(n865), .Q(f33[27]) );
  CFD2QXL \f33_reg[26]  ( .D(s33[26]), .CP(clk), .CD(n865), .Q(f33[26]) );
  CFD2QXL \f33_reg[25]  ( .D(s33[25]), .CP(clk), .CD(n865), .Q(f33[25]) );
  CFD2QXL \f33_reg[24]  ( .D(s33[24]), .CP(clk), .CD(n865), .Q(f33[24]) );
  CFD2QXL \f33_reg[23]  ( .D(s33[23]), .CP(clk), .CD(n865), .Q(f33[23]) );
  CFD2QXL \f33_reg[22]  ( .D(s33[22]), .CP(clk), .CD(n864), .Q(f33[22]) );
  CFD2QXL \f33_reg[21]  ( .D(s33[21]), .CP(clk), .CD(n864), .Q(f33[21]) );
  CFD2QXL \f33_reg[20]  ( .D(s33[20]), .CP(clk), .CD(n864), .Q(f33[20]) );
  CFD2QXL \f41_reg[26]  ( .D(s41[26]), .CP(clk), .CD(n904), .Q(f41[26]) );
  CFD2QXL \f41_reg[25]  ( .D(s41[25]), .CP(clk), .CD(n904), .Q(f41[25]) );
  CFD2QXL \f41_reg[24]  ( .D(s41[24]), .CP(clk), .CD(n904), .Q(f41[24]) );
  CFD2QXL \f41_reg[23]  ( .D(s41[23]), .CP(clk), .CD(n904), .Q(f41[23]) );
  CFD2QXL \f41_reg[22]  ( .D(s41[22]), .CP(clk), .CD(n904), .Q(f41[22]) );
  CFD2QXL \f41_reg[21]  ( .D(s41[21]), .CP(clk), .CD(n904), .Q(f41[21]) );
  CFD2QXL \f41_reg[20]  ( .D(s41[20]), .CP(clk), .CD(n904), .Q(f41[20]) );
  CFD2QXL \f51_reg[18]  ( .D(s51[18]), .CP(clk), .CD(n872), .Q(f51[18]) );
  CFD2QXL \f51_reg[19]  ( .D(s51[19]), .CP(clk), .CD(n872), .Q(f51[19]) );
  CFD2QXL \f51_reg[20]  ( .D(s51[20]), .CP(clk), .CD(n872), .Q(f51[20]) );
  CFD2QXL \f51_reg[21]  ( .D(s51[21]), .CP(clk), .CD(n872), .Q(f51[21]) );
  CFD2QXL \f51_reg[22]  ( .D(s51[22]), .CP(clk), .CD(n872), .Q(f51[22]) );
  CFD2QXL \f51_reg[23]  ( .D(s51[23]), .CP(clk), .CD(n872), .Q(f51[23]) );
  CFD2QXL \f51_reg[24]  ( .D(s51[24]), .CP(clk), .CD(n872), .Q(f51[24]) );
  CFD2QXL \f51_reg[25]  ( .D(s51[25]), .CP(clk), .CD(n872), .Q(f51[25]) );
  CFD2QXL \f51_reg[26]  ( .D(s51[26]), .CP(clk), .CD(n872), .Q(f51[26]) );
  CFD2QXL \f16_reg[26]  ( .D(s16[26]), .CP(clk), .CD(n884), .Q(f16[26]) );
  CFD2QXL \f16_reg[25]  ( .D(s16[25]), .CP(clk), .CD(n884), .Q(f16[25]) );
  CFD2QXL \f16_reg[24]  ( .D(s16[24]), .CP(clk), .CD(n884), .Q(f16[24]) );
  CFD2QXL \f16_reg[23]  ( .D(s16[23]), .CP(clk), .CD(n884), .Q(f16[23]) );
  CFD2QXL \f16_reg[22]  ( .D(s16[22]), .CP(clk), .CD(n884), .Q(f16[22]) );
  CFD2QXL \f16_reg[21]  ( .D(s16[21]), .CP(clk), .CD(n884), .Q(f16[21]) );
  CFD2QXL \f22_reg[27]  ( .D(s22[27]), .CP(clk), .CD(n867), .Q(f22[27]) );
  CFD2QXL \f22_reg[26]  ( .D(s22[26]), .CP(clk), .CD(n867), .Q(f22[26]) );
  CFD2QXL \f22_reg[25]  ( .D(s22[25]), .CP(clk), .CD(n867), .Q(f22[25]) );
  CFD2QXL \f22_reg[24]  ( .D(s22[24]), .CP(clk), .CD(n867), .Q(f22[24]) );
  CFD2QXL \f22_reg[23]  ( .D(s22[23]), .CP(clk), .CD(n867), .Q(f22[23]) );
  CFD2QXL \f22_reg[22]  ( .D(s22[22]), .CP(clk), .CD(n867), .Q(f22[22]) );
  CFD2QXL \f22_reg[21]  ( .D(s22[21]), .CP(clk), .CD(n867), .Q(f22[21]) );
  CFD2QXL \f22_reg[20]  ( .D(s22[20]), .CP(clk), .CD(n867), .Q(f22[20]) );
  CFD2QXL \f27_reg[27]  ( .D(s27[27]), .CP(clk), .CD(n880), .Q(f27[27]) );
  CFD2QXL \f27_reg[26]  ( .D(s27[26]), .CP(clk), .CD(n880), .Q(f27[26]) );
  CFD2QXL \f27_reg[25]  ( .D(s27[25]), .CP(clk), .CD(n879), .Q(f27[25]) );
  CFD2QXL \f27_reg[24]  ( .D(s27[24]), .CP(clk), .CD(n879), .Q(f27[24]) );
  CFD2QXL \f27_reg[23]  ( .D(s27[23]), .CP(clk), .CD(n879), .Q(f27[23]) );
  CFD2QXL \f27_reg[22]  ( .D(s27[22]), .CP(clk), .CD(n879), .Q(f27[22]) );
  CFD2QXL \f27_reg[21]  ( .D(s27[21]), .CP(clk), .CD(n879), .Q(f27[21]) );
  CFD2QXL \f27_reg[20]  ( .D(s27[20]), .CP(clk), .CD(n879), .Q(f27[20]) );
  CFD2QXL \f27_reg[19]  ( .D(s27[19]), .CP(clk), .CD(n879), .Q(f27[19]) );
  CFD2QXL \f34_reg[27]  ( .D(n524), .CP(clk), .CD(n862), .Q(f34[27]) );
  CFD2QXL \f34_reg[26]  ( .D(n522), .CP(clk), .CD(n861), .Q(f34[26]) );
  CFD2QXL \f34_reg[25]  ( .D(n520), .CP(clk), .CD(n861), .Q(f34[25]) );
  CFD2QXL \f34_reg[24]  ( .D(n518), .CP(clk), .CD(n861), .Q(f34[24]) );
  CFD2QXL \f34_reg[23]  ( .D(n516), .CP(clk), .CD(n861), .Q(f34[23]) );
  CFD2QXL \f34_reg[22]  ( .D(n514), .CP(clk), .CD(n860), .Q(f34[22]) );
  CFD2QXL \f34_reg[21]  ( .D(n512), .CP(clk), .CD(n860), .Q(f34[21]) );
  CFD2QXL \f34_reg[20]  ( .D(n510), .CP(clk), .CD(n860), .Q(f34[20]) );
  CFD2QXL \f42_reg[27]  ( .D(n508), .CP(clk), .CD(n877), .Q(f42[27]) );
  CFD2QXL \f42_reg[26]  ( .D(n506), .CP(clk), .CD(n877), .Q(f42[26]) );
  CFD2QXL \f42_reg[25]  ( .D(n504), .CP(clk), .CD(n876), .Q(f42[25]) );
  CFD2QXL \f42_reg[24]  ( .D(n502), .CP(clk), .CD(n876), .Q(f42[24]) );
  CFD2QXL \f42_reg[23]  ( .D(n500), .CP(clk), .CD(n876), .Q(f42[23]) );
  CFD2QXL \f42_reg[22]  ( .D(n498), .CP(clk), .CD(n876), .Q(f42[22]) );
  CFD2QXL \f42_reg[21]  ( .D(n496), .CP(clk), .CD(n876), .Q(f42[21]) );
  CFD2QXL \f42_reg[20]  ( .D(n494), .CP(clk), .CD(n876), .Q(f42[20]) );
  CFD2QXL \f52_reg[27]  ( .D(n492), .CP(clk), .CD(n855), .Q(f52[27]) );
  CFD2QXL \f52_reg[26]  ( .D(n490), .CP(clk), .CD(n854), .Q(f52[26]) );
  CFD2QXL \f52_reg[25]  ( .D(n488), .CP(clk), .CD(n854), .Q(f52[25]) );
  CFD2QXL \f52_reg[24]  ( .D(n486), .CP(clk), .CD(n854), .Q(f52[24]) );
  CFD2QXL \f52_reg[23]  ( .D(n484), .CP(clk), .CD(n854), .Q(f52[23]) );
  CFD2QXL \f52_reg[22]  ( .D(n482), .CP(clk), .CD(n854), .Q(f52[22]) );
  CFD2QXL \f52_reg[21]  ( .D(n480), .CP(clk), .CD(n854), .Q(f52[21]) );
  CFD2QXL \f52_reg[20]  ( .D(n478), .CP(clk), .CD(n854), .Q(f52[20]) );
  CFD2QXL \f52_reg[19]  ( .D(n476), .CP(clk), .CD(n853), .Q(f52[19]) );
  CFD2QXL \f21_reg[31]  ( .D(f11[31]), .CP(clk), .CD(n912), .Q(f21[31]) );
  CFD2QXL \f17_reg[31]  ( .D(s17[31]), .CP(clk), .CD(n882), .Q(f17[31]) );
  CFD2QXL \f01_reg[31]  ( .D(n475), .CP(clk), .CD(n924), .Q(f01[31]) );
  CFD2QXL \f02_reg[31]  ( .D(n474), .CP(clk), .CD(n902), .Q(f02[31]) );
  CFD2QXL \f33_reg[1]  ( .D(s33[1]), .CP(clk), .CD(n863), .Q(f33[1]) );
  CFD2QX1 \f12_reg[25]  ( .D(s12[25]), .CP(clk), .CD(n919), .Q(f12[25]) );
  CFD2QXL \f14_reg[30]  ( .D(s14[30]), .CP(clk), .CD(n895), .Q(f14[30]) );
  CFD2QXL \f30_reg[30]  ( .D(n472), .CP(clk), .CD(n907), .Q(f30[30]) );
  CFD2QXL \f24_reg[19]  ( .D(s24[19]), .CP(clk), .CD(n869), .Q(f24[19]) );
  CFD2QXL \f24_reg[18]  ( .D(s24[18]), .CP(clk), .CD(n869), .Q(f24[18]) );
  CFD2QXL \f24_reg[17]  ( .D(s24[17]), .CP(clk), .CD(n869), .Q(f24[17]) );
  CFD2QXL \f24_reg[16]  ( .D(s24[16]), .CP(clk), .CD(n869), .Q(f24[16]) );
  CFD2QXL \f26_reg[17]  ( .D(s26[17]), .CP(clk), .CD(n891), .Q(f26[17]) );
  CFD2QXL \f26_reg[16]  ( .D(s26[16]), .CP(clk), .CD(n891), .Q(f26[16]) );
  CFD2QXL \f33_reg[19]  ( .D(s33[19]), .CP(clk), .CD(n864), .Q(f33[19]) );
  CFD2QXL \f33_reg[18]  ( .D(s33[18]), .CP(clk), .CD(n864), .Q(f33[18]) );
  CFD2QXL \f33_reg[17]  ( .D(s33[17]), .CP(clk), .CD(n864), .Q(f33[17]) );
  CFD2QXL \f33_reg[16]  ( .D(s33[16]), .CP(clk), .CD(n864), .Q(f33[16]) );
  CFD2QXL \f41_reg[19]  ( .D(s41[19]), .CP(clk), .CD(n904), .Q(f41[19]) );
  CFD2QXL \f41_reg[18]  ( .D(s41[18]), .CP(clk), .CD(n904), .Q(f41[18]) );
  CFD2QXL \f41_reg[17]  ( .D(s41[17]), .CP(clk), .CD(n903), .Q(f41[17]) );
  CFD2QXL \f41_reg[16]  ( .D(s41[16]), .CP(clk), .CD(n903), .Q(f41[16]) );
  CFD2QXL \f51_reg[16]  ( .D(s51[16]), .CP(clk), .CD(n871), .Q(f51[16]) );
  CFD2QXL \f51_reg[17]  ( .D(s51[17]), .CP(clk), .CD(n871), .Q(f51[17]) );
  CFD2QXL \f24_reg[3]  ( .D(s24[3]), .CP(clk), .CD(n868), .Q(f24[3]) );
  CFD2QXL \f33_reg[3]  ( .D(s33[3]), .CP(clk), .CD(n863), .Q(f33[3]) );
  CFD2QXL \f24_reg[1]  ( .D(s24[1]), .CP(clk), .CD(n868), .Q(f24[1]) );
  CFD2QXL \f26_reg[3]  ( .D(s26[3]), .CP(clk), .CD(n890), .Q(f26[3]) );
  CFD2QXL \f26_reg[1]  ( .D(s26[1]), .CP(clk), .CD(n890), .Q(f26[1]) );
  CFD2QXL \f41_reg[3]  ( .D(s41[3]), .CP(clk), .CD(n902), .Q(f41[3]) );
  CFD2QXL \f41_reg[1]  ( .D(s41[1]), .CP(clk), .CD(n902), .Q(f41[1]) );
  CFD2QXL \f51_reg[1]  ( .D(s51[1]), .CP(clk), .CD(n870), .Q(f51[1]) );
  CFD2QXL \f51_reg[3]  ( .D(s51[3]), .CP(clk), .CD(n870), .Q(f51[3]) );
  CFD2QXL \f24_reg[15]  ( .D(s24[15]), .CP(clk), .CD(n869), .Q(f24[15]) );
  CFD2QXL \f24_reg[14]  ( .D(s24[14]), .CP(clk), .CD(n869), .Q(f24[14]) );
  CFD2QXL \f24_reg[13]  ( .D(s24[13]), .CP(clk), .CD(n869), .Q(f24[13]) );
  CFD2QXL \f24_reg[12]  ( .D(s24[12]), .CP(clk), .CD(n869), .Q(f24[12]) );
  CFD2QXL \f24_reg[11]  ( .D(s24[11]), .CP(clk), .CD(n869), .Q(f24[11]) );
  CFD2QXL \f24_reg[10]  ( .D(s24[10]), .CP(clk), .CD(n868), .Q(f24[10]) );
  CFD2QXL \f24_reg[9]  ( .D(s24[9]), .CP(clk), .CD(n868), .Q(f24[9]) );
  CFD2QXL \f24_reg[8]  ( .D(s24[8]), .CP(clk), .CD(n868), .Q(f24[8]) );
  CFD2QXL \f24_reg[7]  ( .D(s24[7]), .CP(clk), .CD(n868), .Q(f24[7]) );
  CFD2QXL \f24_reg[5]  ( .D(s24[5]), .CP(clk), .CD(n868), .Q(f24[5]) );
  CFD2QXL \f24_reg[4]  ( .D(s24[4]), .CP(clk), .CD(n868), .Q(f24[4]) );
  CFD2QXL \f24_reg[0]  ( .D(s24[0]), .CP(clk), .CD(n868), .Q(f24[0]) );
  CFD2QXL \f26_reg[11]  ( .D(s26[11]), .CP(clk), .CD(n891), .Q(f26[11]) );
  CFD2QXL \f26_reg[10]  ( .D(s26[10]), .CP(clk), .CD(n891), .Q(f26[10]) );
  CFD2QXL \f26_reg[9]  ( .D(s26[9]), .CP(clk), .CD(n891), .Q(f26[9]) );
  CFD2QXL \f26_reg[8]  ( .D(s26[8]), .CP(clk), .CD(n890), .Q(f26[8]) );
  CFD2QXL \f26_reg[7]  ( .D(s26[7]), .CP(clk), .CD(n890), .Q(f26[7]) );
  CFD2QXL \f26_reg[5]  ( .D(s26[5]), .CP(clk), .CD(n890), .Q(f26[5]) );
  CFD2QXL \f26_reg[4]  ( .D(s26[4]), .CP(clk), .CD(n890), .Q(f26[4]) );
  CFD2QXL \f26_reg[0]  ( .D(s26[0]), .CP(clk), .CD(n890), .Q(f26[0]) );
  CFD2QXL \f33_reg[15]  ( .D(s33[15]), .CP(clk), .CD(n864), .Q(f33[15]) );
  CFD2QXL \f33_reg[14]  ( .D(s33[14]), .CP(clk), .CD(n864), .Q(f33[14]) );
  CFD2QXL \f33_reg[13]  ( .D(s33[13]), .CP(clk), .CD(n864), .Q(f33[13]) );
  CFD2QXL \f33_reg[12]  ( .D(s33[12]), .CP(clk), .CD(n864), .Q(f33[12]) );
  CFD2QXL \f33_reg[11]  ( .D(s33[11]), .CP(clk), .CD(n864), .Q(f33[11]) );
  CFD2QXL \f33_reg[10]  ( .D(s33[10]), .CP(clk), .CD(n864), .Q(f33[10]) );
  CFD2QXL \f33_reg[9]  ( .D(s33[9]), .CP(clk), .CD(n863), .Q(f33[9]) );
  CFD2QXL \f33_reg[8]  ( .D(s33[8]), .CP(clk), .CD(n863), .Q(f33[8]) );
  CFD2QXL \f33_reg[7]  ( .D(s33[7]), .CP(clk), .CD(n863), .Q(f33[7]) );
  CFD2QXL \f33_reg[5]  ( .D(s33[5]), .CP(clk), .CD(n863), .Q(f33[5]) );
  CFD2QXL \f33_reg[4]  ( .D(s33[4]), .CP(clk), .CD(n863), .Q(f33[4]) );
  CFD2QXL \f33_reg[0]  ( .D(s33[0]), .CP(clk), .CD(n863), .Q(f33[0]) );
  CFD2QXL \f41_reg[11]  ( .D(s41[11]), .CP(clk), .CD(n903), .Q(f41[11]) );
  CFD2QXL \f41_reg[10]  ( .D(s41[10]), .CP(clk), .CD(n903), .Q(f41[10]) );
  CFD2QXL \f41_reg[9]  ( .D(s41[9]), .CP(clk), .CD(n903), .Q(f41[9]) );
  CFD2QXL \f41_reg[8]  ( .D(s41[8]), .CP(clk), .CD(n903), .Q(f41[8]) );
  CFD2QXL \f41_reg[7]  ( .D(s41[7]), .CP(clk), .CD(n903), .Q(f41[7]) );
  CFD2QXL \f41_reg[4]  ( .D(s41[4]), .CP(clk), .CD(n902), .Q(f41[4]) );
  CFD2QXL \f41_reg[0]  ( .D(s41[0]), .CP(clk), .CD(n902), .Q(f41[0]) );
  CFD2QXL \f51_reg[0]  ( .D(s51[0]), .CP(clk), .CD(n870), .Q(f51[0]) );
  CFD2QXL \f51_reg[4]  ( .D(s51[4]), .CP(clk), .CD(n870), .Q(f51[4]) );
  CFD2QXL \f51_reg[5]  ( .D(s51[5]), .CP(clk), .CD(n871), .Q(f51[5]) );
  CFD2QXL \f51_reg[7]  ( .D(s51[7]), .CP(clk), .CD(n871), .Q(f51[7]) );
  CFD2QXL \f51_reg[8]  ( .D(s51[8]), .CP(clk), .CD(n871), .Q(f51[8]) );
  CFD2QXL \f51_reg[9]  ( .D(s51[9]), .CP(clk), .CD(n871), .Q(f51[9]) );
  CFD2QXL \f51_reg[10]  ( .D(s51[10]), .CP(clk), .CD(n871), .Q(f51[10]) );
  CFD2QXL \f51_reg[11]  ( .D(s51[11]), .CP(clk), .CD(n871), .Q(f51[11]) );
  CFD2QXL \f26_reg[15]  ( .D(s26[15]), .CP(clk), .CD(n891), .Q(f26[15]) );
  CFD2QXL \f26_reg[14]  ( .D(s26[14]), .CP(clk), .CD(n891), .Q(f26[14]) );
  CFD2QXL \f26_reg[13]  ( .D(s26[13]), .CP(clk), .CD(n891), .Q(f26[13]) );
  CFD2QXL \f26_reg[12]  ( .D(s26[12]), .CP(clk), .CD(n891), .Q(f26[12]) );
  CFD2QXL \f41_reg[15]  ( .D(s41[15]), .CP(clk), .CD(n903), .Q(f41[15]) );
  CFD2QXL \f41_reg[14]  ( .D(s41[14]), .CP(clk), .CD(n903), .Q(f41[14]) );
  CFD2QXL \f41_reg[13]  ( .D(s41[13]), .CP(clk), .CD(n903), .Q(f41[13]) );
  CFD2QXL \f41_reg[12]  ( .D(s41[12]), .CP(clk), .CD(n903), .Q(f41[12]) );
  CFD2QXL \f51_reg[12]  ( .D(s51[12]), .CP(clk), .CD(n871), .Q(f51[12]) );
  CFD2QXL \f51_reg[13]  ( .D(s51[13]), .CP(clk), .CD(n871), .Q(f51[13]) );
  CFD2QXL \f51_reg[14]  ( .D(s51[14]), .CP(clk), .CD(n871), .Q(f51[14]) );
  CFD2QXL \f51_reg[15]  ( .D(s51[15]), .CP(clk), .CD(n871), .Q(f51[15]) );
  CFD2QXL \f24_reg[6]  ( .D(s24[6]), .CP(clk), .CD(n868), .Q(f24[6]) );
  CFD2QXL \f24_reg[2]  ( .D(s24[2]), .CP(clk), .CD(n868), .Q(f24[2]) );
  CFD2QXL \f26_reg[6]  ( .D(s26[6]), .CP(clk), .CD(n890), .Q(f26[6]) );
  CFD2QXL \f26_reg[2]  ( .D(s26[2]), .CP(clk), .CD(n890), .Q(f26[2]) );
  CFD2QXL \f33_reg[6]  ( .D(s33[6]), .CP(clk), .CD(n863), .Q(f33[6]) );
  CFD2QXL \f33_reg[2]  ( .D(s33[2]), .CP(clk), .CD(n863), .Q(f33[2]) );
  CFD2QXL \f41_reg[6]  ( .D(s41[6]), .CP(clk), .CD(n903), .Q(f41[6]) );
  CFD2QXL \f41_reg[5]  ( .D(s41[5]), .CP(clk), .CD(n903), .Q(f41[5]) );
  CFD2QXL \f41_reg[2]  ( .D(s41[2]), .CP(clk), .CD(n902), .Q(f41[2]) );
  CFD2QXL \f51_reg[2]  ( .D(s51[2]), .CP(clk), .CD(n870), .Q(f51[2]) );
  CFD2QXL \f51_reg[6]  ( .D(s51[6]), .CP(clk), .CD(n871), .Q(f51[6]) );
  CFD2QXL \f14_reg[5]  ( .D(s14[5]), .CP(clk), .CD(n893), .Q(f14[5]) );
  CFD2QXL \f14_reg[9]  ( .D(s14[9]), .CP(clk), .CD(n893), .Q(f14[9]) );
  CFD2QXL \f14_reg[7]  ( .D(s14[7]), .CP(clk), .CD(n893), .Q(f14[7]) );
  CFD2QXL \f30_reg[15]  ( .D(n470), .CP(clk), .CD(n906), .Q(f30[15]) );
  CFD2QXL \f30_reg[12]  ( .D(n468), .CP(clk), .CD(n906), .Q(f30[12]) );
  CFD2QXL \f23_reg[27]  ( .D(s23[27]), .CP(clk), .CD(n914), .Q(f23[27]) );
  CFD2QXL \f30_reg[10]  ( .D(n466), .CP(clk), .CD(n905), .Q(f30[10]) );
  CFD2QXL \f30_reg[11]  ( .D(n465), .CP(clk), .CD(n905), .Q(f30[11]) );
  CFD2QXL \f30_reg[9]  ( .D(n462), .CP(clk), .CD(n905), .Q(f30[9]) );
  CFD2QXL \f30_reg[8]  ( .D(n460), .CP(clk), .CD(n905), .Q(f30[8]) );
  CFD2QXL \f30_reg[6]  ( .D(n458), .CP(clk), .CD(n905), .Q(f30[6]) );
  CFD2QXL \f30_reg[7]  ( .D(n456), .CP(clk), .CD(n905), .Q(f30[7]) );
  CFD2QXL \f30_reg[5]  ( .D(n454), .CP(clk), .CD(n905), .Q(f30[5]) );
  CFD2QXL \f30_reg[4]  ( .D(n452), .CP(clk), .CD(n905), .Q(f30[4]) );
  CFD2QXL \f30_reg[3]  ( .D(n450), .CP(clk), .CD(n905), .Q(f30[3]) );
  CFD2QXL \f30_reg[2]  ( .D(n448), .CP(clk), .CD(n905), .Q(f30[2]) );
  CFD2QXL \f31_reg[27]  ( .D(s31[27]), .CP(clk), .CD(n909), .Q(f31[27]) );
  CFD2QXL \f14_reg[15]  ( .D(s14[15]), .CP(clk), .CD(n893), .Q(f14[15]) );
  CFD2QXL \f03_reg[30]  ( .D(n446), .CP(clk), .CD(n890), .Q(f03[30]) );
  CFD2QXL \f16_reg[20]  ( .D(s16[20]), .CP(clk), .CD(n884), .Q(f16[20]) );
  CFD2QXL \f16_reg[19]  ( .D(s16[19]), .CP(clk), .CD(n884), .Q(f16[19]) );
  CFD2QXL \f16_reg[18]  ( .D(s16[18]), .CP(clk), .CD(n884), .Q(f16[18]) );
  CFD2QXL \f16_reg[17]  ( .D(s16[17]), .CP(clk), .CD(n884), .Q(f16[17]) );
  CFD2QXL \f16_reg[16]  ( .D(s16[16]), .CP(clk), .CD(n884), .Q(f16[16]) );
  CFD2QXL \f22_reg[19]  ( .D(s22[19]), .CP(clk), .CD(n867), .Q(f22[19]) );
  CFD2QXL \f22_reg[18]  ( .D(s22[18]), .CP(clk), .CD(n867), .Q(f22[18]) );
  CFD2QXL \f22_reg[17]  ( .D(s22[17]), .CP(clk), .CD(n867), .Q(f22[17]) );
  CFD2QXL \f22_reg[16]  ( .D(s22[16]), .CP(clk), .CD(n866), .Q(f22[16]) );
  CFD2QXL \f27_reg[18]  ( .D(s27[18]), .CP(clk), .CD(n879), .Q(f27[18]) );
  CFD2QXL \f27_reg[17]  ( .D(s27[17]), .CP(clk), .CD(n879), .Q(f27[17]) );
  CFD2QXL \f27_reg[16]  ( .D(s27[16]), .CP(clk), .CD(n879), .Q(f27[16]) );
  CFD2QXL \f34_reg[19]  ( .D(n444), .CP(clk), .CD(n860), .Q(f34[19]) );
  CFD2QXL \f34_reg[18]  ( .D(n442), .CP(clk), .CD(n860), .Q(f34[18]) );
  CFD2QXL \f34_reg[17]  ( .D(n440), .CP(clk), .CD(n859), .Q(f34[17]) );
  CFD2QXL \f34_reg[16]  ( .D(n438), .CP(clk), .CD(n859), .Q(f34[16]) );
  CFD2QXL \f42_reg[19]  ( .D(n436), .CP(clk), .CD(n876), .Q(f42[19]) );
  CFD2QXL \f42_reg[18]  ( .D(n434), .CP(clk), .CD(n875), .Q(f42[18]) );
  CFD2QXL \f42_reg[17]  ( .D(n432), .CP(clk), .CD(n875), .Q(f42[17]) );
  CFD2QXL \f42_reg[16]  ( .D(n430), .CP(clk), .CD(n875), .Q(f42[16]) );
  CFD2QXL \f52_reg[18]  ( .D(n428), .CP(clk), .CD(n853), .Q(f52[18]) );
  CFD2QXL \f52_reg[17]  ( .D(n426), .CP(clk), .CD(n853), .Q(f52[17]) );
  CFD2QXL \f52_reg[16]  ( .D(n424), .CP(clk), .CD(n853), .Q(f52[16]) );
  CFD2QXL \f22_reg[3]  ( .D(s22[3]), .CP(clk), .CD(n865), .Q(f22[3]) );
  CFD2QXL \f34_reg[3]  ( .D(n422), .CP(clk), .CD(n856), .Q(f34[3]) );
  CFD2QXL \f16_reg[3]  ( .D(s16[3]), .CP(clk), .CD(n883), .Q(f16[3]) );
  CFD2QXL \f16_reg[1]  ( .D(s16[1]), .CP(clk), .CD(n883), .Q(f16[1]) );
  CFD2QXL \f22_reg[1]  ( .D(s22[1]), .CP(clk), .CD(n865), .Q(f22[1]) );
  CFD2QXL \f27_reg[3]  ( .D(s27[3]), .CP(clk), .CD(n878), .Q(f27[3]) );
  CFD2QXL \f27_reg[1]  ( .D(s27[1]), .CP(clk), .CD(n878), .Q(f27[1]) );
  CFD2QXL \f42_reg[3]  ( .D(n420), .CP(clk), .CD(n873), .Q(f42[3]) );
  CFD2QXL \f42_reg[1]  ( .D(n418), .CP(clk), .CD(n873), .Q(f42[1]) );
  CFD2QXL \f52_reg[3]  ( .D(n416), .CP(clk), .CD(n851), .Q(f52[3]) );
  CFD2QXL \f52_reg[1]  ( .D(n414), .CP(clk), .CD(n851), .Q(f52[1]) );
  CFD2QXL \f16_reg[11]  ( .D(s16[11]), .CP(clk), .CD(n883), .Q(f16[11]) );
  CFD2QXL \f16_reg[10]  ( .D(s16[10]), .CP(clk), .CD(n883), .Q(f16[10]) );
  CFD2QXL \f16_reg[9]  ( .D(s16[9]), .CP(clk), .CD(n883), .Q(f16[9]) );
  CFD2QXL \f16_reg[8]  ( .D(s16[8]), .CP(clk), .CD(n883), .Q(f16[8]) );
  CFD2QXL \f16_reg[7]  ( .D(s16[7]), .CP(clk), .CD(n883), .Q(f16[7]) );
  CFD2QXL \f16_reg[4]  ( .D(s16[4]), .CP(clk), .CD(n883), .Q(f16[4]) );
  CFD2QXL \f16_reg[0]  ( .D(s16[0]), .CP(clk), .CD(n882), .Q(f16[0]) );
  CFD2QXL \f22_reg[15]  ( .D(s22[15]), .CP(clk), .CD(n866), .Q(f22[15]) );
  CFD2QXL \f22_reg[14]  ( .D(s22[14]), .CP(clk), .CD(n866), .Q(f22[14]) );
  CFD2QXL \f22_reg[13]  ( .D(s22[13]), .CP(clk), .CD(n866), .Q(f22[13]) );
  CFD2QXL \f22_reg[12]  ( .D(s22[12]), .CP(clk), .CD(n866), .Q(f22[12]) );
  CFD2QXL \f22_reg[11]  ( .D(s22[11]), .CP(clk), .CD(n866), .Q(f22[11]) );
  CFD2QXL \f22_reg[10]  ( .D(s22[10]), .CP(clk), .CD(n866), .Q(f22[10]) );
  CFD2QXL \f22_reg[9]  ( .D(s22[9]), .CP(clk), .CD(n866), .Q(f22[9]) );
  CFD2QXL \f22_reg[8]  ( .D(s22[8]), .CP(clk), .CD(n866), .Q(f22[8]) );
  CFD2QXL \f22_reg[7]  ( .D(s22[7]), .CP(clk), .CD(n866), .Q(f22[7]) );
  CFD2QXL \f22_reg[5]  ( .D(s22[5]), .CP(clk), .CD(n866), .Q(f22[5]) );
  CFD2QXL \f22_reg[4]  ( .D(s22[4]), .CP(clk), .CD(n866), .Q(f22[4]) );
  CFD2QXL \f22_reg[0]  ( .D(s22[0]), .CP(clk), .CD(n865), .Q(f22[0]) );
  CFD2QXL \f27_reg[11]  ( .D(s27[11]), .CP(clk), .CD(n878), .Q(f27[11]) );
  CFD2QXL \f27_reg[10]  ( .D(s27[10]), .CP(clk), .CD(n878), .Q(f27[10]) );
  CFD2QXL \f27_reg[9]  ( .D(s27[9]), .CP(clk), .CD(n878), .Q(f27[9]) );
  CFD2QXL \f27_reg[8]  ( .D(s27[8]), .CP(clk), .CD(n878), .Q(f27[8]) );
  CFD2QXL \f27_reg[7]  ( .D(s27[7]), .CP(clk), .CD(n878), .Q(f27[7]) );
  CFD2QXL \f27_reg[5]  ( .D(s27[5]), .CP(clk), .CD(n878), .Q(f27[5]) );
  CFD2QXL \f27_reg[4]  ( .D(s27[4]), .CP(clk), .CD(n878), .Q(f27[4]) );
  CFD2QXL \f27_reg[0]  ( .D(s27[0]), .CP(clk), .CD(n878), .Q(f27[0]) );
  CFD2QXL \f34_reg[15]  ( .D(n412), .CP(clk), .CD(n859), .Q(f34[15]) );
  CFD2QXL \f34_reg[14]  ( .D(n410), .CP(clk), .CD(n859), .Q(f34[14]) );
  CFD2QXL \f34_reg[13]  ( .D(n408), .CP(clk), .CD(n858), .Q(f34[13]) );
  CFD2QXL \f34_reg[12]  ( .D(n406), .CP(clk), .CD(n858), .Q(f34[12]) );
  CFD2QXL \f34_reg[11]  ( .D(n404), .CP(clk), .CD(n858), .Q(f34[11]) );
  CFD2QXL \f34_reg[10]  ( .D(n402), .CP(clk), .CD(n858), .Q(f34[10]) );
  CFD2QXL \f34_reg[9]  ( .D(n400), .CP(clk), .CD(n857), .Q(f34[9]) );
  CFD2QXL \f34_reg[8]  ( .D(n398), .CP(clk), .CD(n857), .Q(f34[8]) );
  CFD2QXL \f34_reg[7]  ( .D(n396), .CP(clk), .CD(n857), .Q(f34[7]) );
  CFD2QXL \f34_reg[5]  ( .D(n394), .CP(clk), .CD(n857), .Q(f34[5]) );
  CFD2QXL \f34_reg[4]  ( .D(n392), .CP(clk), .CD(n856), .Q(f34[4]) );
  CFD2QXL \f34_reg[0]  ( .D(n390), .CP(clk), .CD(n855), .Q(f34[0]) );
  CFD2QXL \f42_reg[11]  ( .D(n388), .CP(clk), .CD(n874), .Q(f42[11]) );
  CFD2QXL \f42_reg[10]  ( .D(n386), .CP(clk), .CD(n874), .Q(f42[10]) );
  CFD2QXL \f42_reg[9]  ( .D(n384), .CP(clk), .CD(n874), .Q(f42[9]) );
  CFD2QXL \f42_reg[8]  ( .D(n382), .CP(clk), .CD(n874), .Q(f42[8]) );
  CFD2QXL \f42_reg[7]  ( .D(n380), .CP(clk), .CD(n874), .Q(f42[7]) );
  CFD2QXL \f42_reg[4]  ( .D(n378), .CP(clk), .CD(n873), .Q(f42[4]) );
  CFD2QXL \f42_reg[0]  ( .D(n376), .CP(clk), .CD(n873), .Q(f42[0]) );
  CFD2QXL \f52_reg[11]  ( .D(n374), .CP(clk), .CD(n852), .Q(f52[11]) );
  CFD2QXL \f52_reg[10]  ( .D(n372), .CP(clk), .CD(n852), .Q(f52[10]) );
  CFD2QXL \f52_reg[9]  ( .D(n370), .CP(clk), .CD(n852), .Q(f52[9]) );
  CFD2QXL \f52_reg[8]  ( .D(n368), .CP(clk), .CD(n852), .Q(f52[8]) );
  CFD2QXL \f52_reg[7]  ( .D(n366), .CP(clk), .CD(n852), .Q(f52[7]) );
  CFD2QXL \f52_reg[5]  ( .D(n364), .CP(clk), .CD(n851), .Q(f52[5]) );
  CFD2QXL \f52_reg[4]  ( .D(n362), .CP(clk), .CD(n851), .Q(f52[4]) );
  CFD2QXL \f52_reg[0]  ( .D(n360), .CP(clk), .CD(n850), .Q(f52[0]) );
  CFD2QXL \f16_reg[14]  ( .D(s16[14]), .CP(clk), .CD(n884), .Q(f16[14]) );
  CFD2QXL \f16_reg[13]  ( .D(s16[13]), .CP(clk), .CD(n883), .Q(f16[13]) );
  CFD2QXL \f16_reg[12]  ( .D(s16[12]), .CP(clk), .CD(n883), .Q(f16[12]) );
  CFD2QXL \f27_reg[15]  ( .D(s27[15]), .CP(clk), .CD(n879), .Q(f27[15]) );
  CFD2QXL \f27_reg[14]  ( .D(s27[14]), .CP(clk), .CD(n879), .Q(f27[14]) );
  CFD2QXL \f27_reg[13]  ( .D(s27[13]), .CP(clk), .CD(n879), .Q(f27[13]) );
  CFD2QXL \f27_reg[12]  ( .D(s27[12]), .CP(clk), .CD(n878), .Q(f27[12]) );
  CFD2QXL \f42_reg[15]  ( .D(n358), .CP(clk), .CD(n875), .Q(f42[15]) );
  CFD2QXL \f42_reg[14]  ( .D(n356), .CP(clk), .CD(n875), .Q(f42[14]) );
  CFD2QXL \f42_reg[13]  ( .D(n354), .CP(clk), .CD(n875), .Q(f42[13]) );
  CFD2QXL \f42_reg[12]  ( .D(n352), .CP(clk), .CD(n874), .Q(f42[12]) );
  CFD2QXL \f52_reg[15]  ( .D(n350), .CP(clk), .CD(n853), .Q(f52[15]) );
  CFD2QXL \f52_reg[14]  ( .D(n348), .CP(clk), .CD(n853), .Q(f52[14]) );
  CFD2QXL \f52_reg[13]  ( .D(n346), .CP(clk), .CD(n852), .Q(f52[13]) );
  CFD2QXL \f52_reg[12]  ( .D(n344), .CP(clk), .CD(n852), .Q(f52[12]) );
  CFD2QXL \f16_reg[6]  ( .D(s16[6]), .CP(clk), .CD(n883), .Q(f16[6]) );
  CFD2QXL \f16_reg[5]  ( .D(s16[5]), .CP(clk), .CD(n883), .Q(f16[5]) );
  CFD2QXL \f16_reg[2]  ( .D(s16[2]), .CP(clk), .CD(n883), .Q(f16[2]) );
  CFD2QXL \f22_reg[6]  ( .D(s22[6]), .CP(clk), .CD(n866), .Q(f22[6]) );
  CFD2QXL \f22_reg[2]  ( .D(s22[2]), .CP(clk), .CD(n865), .Q(f22[2]) );
  CFD2QXL \f27_reg[6]  ( .D(s27[6]), .CP(clk), .CD(n878), .Q(f27[6]) );
  CFD2QXL \f27_reg[2]  ( .D(s27[2]), .CP(clk), .CD(n878), .Q(f27[2]) );
  CFD2QXL \f34_reg[6]  ( .D(n342), .CP(clk), .CD(n857), .Q(f34[6]) );
  CFD2QXL \f34_reg[2]  ( .D(n340), .CP(clk), .CD(n856), .Q(f34[2]) );
  CFD2QXL \f42_reg[6]  ( .D(n338), .CP(clk), .CD(n874), .Q(f42[6]) );
  CFD2QXL \f42_reg[5]  ( .D(n336), .CP(clk), .CD(n873), .Q(f42[5]) );
  CFD2QXL \f42_reg[2]  ( .D(n334), .CP(clk), .CD(n873), .Q(f42[2]) );
  CFD2QXL \f52_reg[6]  ( .D(n332), .CP(clk), .CD(n851), .Q(f52[6]) );
  CFD2QXL \f52_reg[2]  ( .D(n330), .CP(clk), .CD(n851), .Q(f52[2]) );
  CFD2QXL \f21_reg[30]  ( .D(n329), .CP(clk), .CD(n912), .Q(f21[30]) );
  CFD2QXL \f21_reg[4]  ( .D(n326), .CP(clk), .CD(n910), .Q(f21[4]) );
  CFD2QXL \f21_reg[2]  ( .D(n325), .CP(clk), .CD(n910), .Q(f21[2]) );
  CFD2QXL \f21_reg[14]  ( .D(n323), .CP(clk), .CD(n911), .Q(f21[14]) );
  CFD2QXL \f21_reg[12]  ( .D(n322), .CP(clk), .CD(n910), .Q(f21[12]) );
  CFD2QXL \f21_reg[9]  ( .D(n319), .CP(clk), .CD(n910), .Q(f21[9]) );
  CFD2QXL \f21_reg[5]  ( .D(n316), .CP(clk), .CD(n910), .Q(f21[5]) );
  CFD2QXL \f17_reg[30]  ( .D(s17[30]), .CP(clk), .CD(n882), .Q(f17[30]) );
  CFD2QXL \f16_reg[15]  ( .D(s16[15]), .CP(clk), .CD(n884), .Q(f16[15]) );
  CFD2QXL \f17_reg[29]  ( .D(s17[29]), .CP(clk), .CD(n882), .Q(f17[29]) );
  CFD2QXL \f03_reg[28]  ( .D(n315), .CP(clk), .CD(n889), .Q(f03[28]) );
  CFD2QXL \f14_reg[29]  ( .D(s14[29]), .CP(clk), .CD(n895), .Q(f14[29]) );
  CFD2QXL \f14_reg[28]  ( .D(s14[28]), .CP(clk), .CD(n894), .Q(f14[28]) );
  CFD2QXL \f30_reg[29]  ( .D(n314), .CP(clk), .CD(n907), .Q(f30[29]) );
  CFD2QXL \f30_reg[28]  ( .D(n313), .CP(clk), .CD(n907), .Q(f30[28]) );
  CFD2QXL \f23_reg[30]  ( .D(s23[30]), .CP(clk), .CD(n914), .Q(f23[30]) );
  CFD2QXL \f23_reg[28]  ( .D(s23[28]), .CP(clk), .CD(n914), .Q(f23[28]) );
  CFD2QXL \f31_reg[30]  ( .D(s31[30]), .CP(clk), .CD(n909), .Q(f31[30]) );
  CFD2QXL \f31_reg[28]  ( .D(s31[28]), .CP(clk), .CD(n909), .Q(f31[28]) );
  CFD2QXL \f31_reg[26]  ( .D(s31[26]), .CP(clk), .CD(n909), .Q(f31[26]) );
  CFD2QXL \f23_reg[26]  ( .D(s23[26]), .CP(clk), .CD(n914), .Q(f23[26]) );
  CFD2QXL \f21_reg[29]  ( .D(f11[29]), .CP(clk), .CD(n912), .Q(f21[29]) );
  CFD2QXL \f21_reg[28]  ( .D(n312), .CP(clk), .CD(n912), .Q(f21[28]) );
  CFD2QXL \f14_reg[26]  ( .D(s14[26]), .CP(clk), .CD(n894), .Q(f14[26]) );
  CFD2QXL \f13_reg[30]  ( .D(n311), .CP(clk), .CD(n902), .Q(f13[30]) );
  CFD2QXL \f17_reg[28]  ( .D(s17[28]), .CP(clk), .CD(n882), .Q(f17[28]) );
  CFD2QXL \f14_reg[25]  ( .D(s14[25]), .CP(clk), .CD(n894), .Q(f14[25]) );
  CFD2QXL \f14_reg[24]  ( .D(s14[24]), .CP(clk), .CD(n894), .Q(f14[24]) );
  CFD2QXL \f21_reg[7]  ( .D(n309), .CP(clk), .CD(n910), .Q(f21[7]) );
  CFD2QXL \f21_reg[11]  ( .D(n306), .CP(clk), .CD(n910), .Q(f21[11]) );
  CFD2QXL \f01_reg[30]  ( .D(n305), .CP(clk), .CD(n924), .Q(f01[30]) );
  CFD2QXL \f01_reg[28]  ( .D(n304), .CP(clk), .CD(n924), .Q(f01[28]) );
  CFD2QXL \f02_reg[30]  ( .D(n303), .CP(clk), .CD(n902), .Q(f02[30]) );
  CFD2QXL \f02_reg[28]  ( .D(n302), .CP(clk), .CD(n901), .Q(f02[28]) );
  CFD2QXL \f11_reg[30]  ( .D(n301), .CP(clk), .CD(n917), .Q(f11[30]) );
  CFD2QXL \f14_reg[22]  ( .D(s14[22]), .CP(clk), .CD(n894), .Q(f14[22]) );
  CFD2QXL \f14_reg[27]  ( .D(s14[27]), .CP(clk), .CD(n894), .Q(f14[27]) );
  CFD2QXL \f30_reg[27]  ( .D(n300), .CP(clk), .CD(n907), .Q(f30[27]) );
  CFD2QXL \f30_reg[26]  ( .D(n299), .CP(clk), .CD(n907), .Q(f30[26]) );
  CFD2QXL \f11_reg[28]  ( .D(n298), .CP(clk), .CD(n917), .Q(f11[28]) );
  CFD2QXL \f03_reg[29]  ( .D(n297), .CP(clk), .CD(n889), .Q(f03[29]) );
  CFD2QXL \f21_reg[27]  ( .D(n296), .CP(clk), .CD(n912), .Q(f21[27]) );
  CFD2QXL \f21_reg[26]  ( .D(n294), .CP(clk), .CD(n912), .Q(f21[26]) );
  CFD2QXL \f30_reg[24]  ( .D(f21[24]), .CP(clk), .CD(n906), .Q(f30[24]) );
  CFD2QXL \f17_reg[27]  ( .D(s17[27]), .CP(clk), .CD(n882), .Q(f17[27]) );
  CFD2QXL \f14_reg[21]  ( .D(s14[21]), .CP(clk), .CD(n894), .Q(f14[21]) );
  CFD2QXL \f11_reg[31]  ( .D(f01[31]), .CP(clk), .CD(n917), .Q(f11[31]) );
  CFD2QXL \f21_reg[25]  ( .D(n293), .CP(clk), .CD(n911), .Q(f21[25]) );
  CFD2QXL \f21_reg[24]  ( .D(n290), .CP(clk), .CD(n911), .Q(f21[24]) );
  CFD2QXL \f30_reg[23]  ( .D(n289), .CP(clk), .CD(n906), .Q(f30[23]) );
  CFD2QXL \f17_reg[26]  ( .D(s17[26]), .CP(clk), .CD(n882), .Q(f17[26]) );
  CFD2QXL \f21_reg[20]  ( .D(n288), .CP(clk), .CD(n911), .Q(f21[20]) );
  CFD2QXL \f21_reg[23]  ( .D(n286), .CP(clk), .CD(n911), .Q(f21[23]) );
  CFD2QXL \f14_reg[23]  ( .D(s14[23]), .CP(clk), .CD(n894), .Q(f14[23]) );
  CFD2QXL \f30_reg[22]  ( .D(f21[22]), .CP(clk), .CD(n906), .Q(f30[22]) );
  CFD2QXL \f23_reg[31]  ( .D(s23[31]), .CP(clk), .CD(n914), .Q(f23[31]) );
  CFD2QXL \f17_reg[25]  ( .D(s17[25]), .CP(clk), .CD(n882), .Q(f17[25]) );
  CFD2QXL \f03_reg[27]  ( .D(n285), .CP(clk), .CD(n889), .Q(f03[27]) );
  CFD2QXL \f17_reg[21]  ( .D(s17[21]), .CP(clk), .CD(n882), .Q(f17[21]) );
  CFD2QXL \f30_reg[25]  ( .D(f21[25]), .CP(clk), .CD(n907), .Q(f30[25]) );
  CFD2QXL \f21_reg[22]  ( .D(n284), .CP(clk), .CD(n911), .Q(f21[22]) );
  CFD2QXL \f12_reg[30]  ( .D(s12[30]), .CP(clk), .CD(n919), .Q(f12[30]) );
  CFD2QXL \f17_reg[22]  ( .D(s17[22]), .CP(clk), .CD(n882), .Q(f17[22]) );
  CFD2QXL \f17_reg[24]  ( .D(s17[24]), .CP(clk), .CD(n882), .Q(f17[24]) );
  CFD2QXL \f17_reg[20]  ( .D(s17[20]), .CP(clk), .CD(n882), .Q(f17[20]) );
  CFD2QXL \f13_reg[31]  ( .D(f02[31]), .CP(clk), .CD(n902), .Q(f13[31]) );
  CFD2QXL \f17_reg[23]  ( .D(s17[23]), .CP(clk), .CD(n882), .Q(f17[23]) );
  CFD2QXL \f12_reg[31]  ( .D(s12[31]), .CP(clk), .CD(n919), .Q(f12[31]) );
  CFD2QX1 \f03_reg[13]  ( .D(n282), .CP(clk), .CD(n887), .Q(f03[13]) );
  CFD2QXL \f23_reg[29]  ( .D(s23[29]), .CP(clk), .CD(n914), .Q(f23[29]) );
  CFD2QXL \f30_reg[21]  ( .D(n280), .CP(clk), .CD(n906), .Q(f30[21]) );
  CFD2QXL \f15_reg[2]  ( .D(s15[2]), .CP(clk), .CD(n856), .Q(f15[2]) );
  CFD2QXL \f32_reg[31]  ( .D(s32[31]), .CP(clk), .CD(n877), .Q(f32[31]) );
  CFD2QXL \f32_reg[30]  ( .D(s32[30]), .CP(clk), .CD(n877), .Q(f32[30]) );
  CFD2QXL \f32_reg[29]  ( .D(s32[29]), .CP(clk), .CD(n877), .Q(f32[29]) );
  CFD2QXL \f32_reg[28]  ( .D(s32[28]), .CP(clk), .CD(n877), .Q(f32[28]) );
  CFD2QXL \f32_reg[0]  ( .D(s32[0]), .CP(clk), .CD(n873), .Q(f32[0]) );
  CFD2QXL \f43_reg[31]  ( .D(s43[31]), .CP(clk), .CD(n855), .Q(f43[31]) );
  CFD2QXL \f43_reg[30]  ( .D(s43[30]), .CP(clk), .CD(n855), .Q(f43[30]) );
  CFD2QXL \f43_reg[29]  ( .D(s43[29]), .CP(clk), .CD(n855), .Q(f43[29]) );
  CFD2QXL \f43_reg[28]  ( .D(s43[28]), .CP(clk), .CD(n855), .Q(f43[28]) );
  CFD2QXL \f43_reg[1]  ( .D(s43[1]), .CP(clk), .CD(n851), .Q(f43[1]) );
  CFD2QXL \f43_reg[0]  ( .D(s43[0]), .CP(clk), .CD(n851), .Q(f43[0]) );
  CFD2QXL \res_d_reg[0]  ( .D(res_temp[0]), .CP(clk), .CD(n850), .Q(res_d[0])
         );
  CFD2QXL \res_d_reg[28]  ( .D(res_temp[28]), .CP(clk), .CD(n846), .Q(
        res_d[28]) );
  CFD2QXL \res_d_reg[29]  ( .D(res_temp[29]), .CP(clk), .CD(n846), .Q(
        res_d[29]) );
  CFD2QXL \res_d_reg[30]  ( .D(res_temp[30]), .CP(clk), .CD(n846), .Q(
        res_d[30]) );
  CFD2QXL \res_d_reg[31]  ( .D(res_temp[31]), .CP(clk), .CD(n846), .Q(
        res_d[31]) );
  CFD2QXL all_in_reg ( .D(N6), .CP(clk), .CD(n924), .Q(all_in) );
  CFD2QXL all_in1_reg ( .D(n278), .CP(clk), .CD(n924), .Q(all_in1) );
  CFD2QXL all_in2_reg ( .D(n276), .CP(clk), .CD(n925), .Q(all_in2) );
  CFD2QXL all_in3_reg ( .D(n274), .CP(clk), .CD(n925), .Q(all_in3) );
  CFD2QXL all_in4_reg ( .D(n272), .CP(clk), .CD(n925), .Q(all_in4) );
  CFD2QXL all_in5_reg ( .D(n270), .CP(clk), .CD(n925), .Q(all_in5) );
  CFD2QXL all_in6_reg ( .D(n268), .CP(clk), .CD(n925), .Q(all_in6) );
  CFD2QXL all_in7_reg ( .D(n266), .CP(clk), .CD(n925), .Q(all_in7) );
  CFD2QXL \f15_reg[31]  ( .D(s15[31]), .CP(clk), .CD(n863), .Q(f15[31]) );
  CFD2QXL \f15_reg[30]  ( .D(s15[30]), .CP(clk), .CD(n862), .Q(f15[30]) );
  CFD2QXL \f15_reg[29]  ( .D(s15[29]), .CP(clk), .CD(n862), .Q(f15[29]) );
  CFD2QXL \f15_reg[28]  ( .D(s15[28]), .CP(clk), .CD(n862), .Q(f15[28]) );
  CFD2QXL \f15_reg[26]  ( .D(s15[26]), .CP(clk), .CD(n862), .Q(f15[26]) );
  CFD2QXL \f15_reg[25]  ( .D(s15[25]), .CP(clk), .CD(n861), .Q(f15[25]) );
  CFD2QXL \f15_reg[24]  ( .D(s15[24]), .CP(clk), .CD(n861), .Q(f15[24]) );
  CFD2QXL \f15_reg[23]  ( .D(s15[23]), .CP(clk), .CD(n861), .Q(f15[23]) );
  CFD2QXL \f15_reg[22]  ( .D(s15[22]), .CP(clk), .CD(n861), .Q(f15[22]) );
  CFD2QXL \f15_reg[21]  ( .D(s15[21]), .CP(clk), .CD(n860), .Q(f15[21]) );
  CFD2QXL \f15_reg[20]  ( .D(s15[20]), .CP(clk), .CD(n860), .Q(f15[20]) );
  CFD2QXL \f15_reg[19]  ( .D(s15[19]), .CP(clk), .CD(n860), .Q(f15[19]) );
  CFD2QXL \f15_reg[18]  ( .D(s15[18]), .CP(clk), .CD(n860), .Q(f15[18]) );
  CFD2QXL \f15_reg[17]  ( .D(s15[17]), .CP(clk), .CD(n859), .Q(f15[17]) );
  CFD2QXL \f15_reg[16]  ( .D(s15[16]), .CP(clk), .CD(n859), .Q(f15[16]) );
  CFD2QXL \f15_reg[15]  ( .D(s15[15]), .CP(clk), .CD(n859), .Q(f15[15]) );
  CFD2QXL \f15_reg[14]  ( .D(s15[14]), .CP(clk), .CD(n859), .Q(f15[14]) );
  CFD2QXL \f15_reg[13]  ( .D(s15[13]), .CP(clk), .CD(n859), .Q(f15[13]) );
  CFD2QXL \f15_reg[12]  ( .D(s15[12]), .CP(clk), .CD(n858), .Q(f15[12]) );
  CFD2QXL \f15_reg[11]  ( .D(s15[11]), .CP(clk), .CD(n858), .Q(f15[11]) );
  CFD2QXL \f15_reg[10]  ( .D(s15[10]), .CP(clk), .CD(n858), .Q(f15[10]) );
  CFD2QXL \f15_reg[9]  ( .D(s15[9]), .CP(clk), .CD(n858), .Q(f15[9]) );
  CFD2QXL \f15_reg[8]  ( .D(s15[8]), .CP(clk), .CD(n857), .Q(f15[8]) );
  CFD2QXL \f15_reg[7]  ( .D(s15[7]), .CP(clk), .CD(n857), .Q(f15[7]) );
  CFD2QXL \f15_reg[6]  ( .D(s15[6]), .CP(clk), .CD(n857), .Q(f15[6]) );
  CFD2QXL \f15_reg[5]  ( .D(s15[5]), .CP(clk), .CD(n857), .Q(f15[5]) );
  CFD2QXL \f15_reg[4]  ( .D(s15[4]), .CP(clk), .CD(n856), .Q(f15[4]) );
  CFD2QXL \f15_reg[3]  ( .D(s15[3]), .CP(clk), .CD(n856), .Q(f15[3]) );
  CFD2QXL \f15_reg[0]  ( .D(s15[0]), .CP(clk), .CD(n856), .Q(f15[0]) );
  CFD2QXL \f25_reg[31]  ( .D(n262), .CP(clk), .CD(n863), .Q(f25[31]) );
  CFD2QXL \f25_reg[30]  ( .D(n260), .CP(clk), .CD(n862), .Q(f25[30]) );
  CFD2QXL \f25_reg[29]  ( .D(n258), .CP(clk), .CD(n862), .Q(f25[29]) );
  CFD2QXL \f25_reg[28]  ( .D(n256), .CP(clk), .CD(n862), .Q(f25[28]) );
  CFD2QXL \f25_reg[27]  ( .D(n254), .CP(clk), .CD(n862), .Q(f25[27]) );
  CFD2QXL \f25_reg[26]  ( .D(n252), .CP(clk), .CD(n861), .Q(f25[26]) );
  CFD2QXL \f25_reg[25]  ( .D(n250), .CP(clk), .CD(n861), .Q(f25[25]) );
  CFD2QXL \f25_reg[24]  ( .D(n248), .CP(clk), .CD(n861), .Q(f25[24]) );
  CFD2QXL \f25_reg[23]  ( .D(n246), .CP(clk), .CD(n861), .Q(f25[23]) );
  CFD2QXL \f25_reg[22]  ( .D(n244), .CP(clk), .CD(n861), .Q(f25[22]) );
  CFD2QXL \f25_reg[21]  ( .D(n242), .CP(clk), .CD(n860), .Q(f25[21]) );
  CFD2QXL \f25_reg[20]  ( .D(n240), .CP(clk), .CD(n860), .Q(f25[20]) );
  CFD2QXL \f25_reg[19]  ( .D(n238), .CP(clk), .CD(n860), .Q(f25[19]) );
  CFD2QXL \f25_reg[18]  ( .D(n236), .CP(clk), .CD(n860), .Q(f25[18]) );
  CFD2QXL \f25_reg[17]  ( .D(n234), .CP(clk), .CD(n859), .Q(f25[17]) );
  CFD2QXL \f25_reg[16]  ( .D(n232), .CP(clk), .CD(n859), .Q(f25[16]) );
  CFD2QXL \f25_reg[15]  ( .D(n230), .CP(clk), .CD(n859), .Q(f25[15]) );
  CFD2QXL \f25_reg[14]  ( .D(n228), .CP(clk), .CD(n859), .Q(f25[14]) );
  CFD2QXL \f25_reg[13]  ( .D(n226), .CP(clk), .CD(n858), .Q(f25[13]) );
  CFD2QXL \f25_reg[12]  ( .D(n224), .CP(clk), .CD(n858), .Q(f25[12]) );
  CFD2QXL \f25_reg[11]  ( .D(n222), .CP(clk), .CD(n858), .Q(f25[11]) );
  CFD2QXL \f25_reg[10]  ( .D(n220), .CP(clk), .CD(n858), .Q(f25[10]) );
  CFD2QXL \f25_reg[9]  ( .D(n218), .CP(clk), .CD(n858), .Q(f25[9]) );
  CFD2QXL \f25_reg[8]  ( .D(n216), .CP(clk), .CD(n857), .Q(f25[8]) );
  CFD2QXL \f25_reg[7]  ( .D(n214), .CP(clk), .CD(n857), .Q(f25[7]) );
  CFD2QXL \f25_reg[6]  ( .D(n212), .CP(clk), .CD(n857), .Q(f25[6]) );
  CFD2QXL \f25_reg[5]  ( .D(n210), .CP(clk), .CD(n857), .Q(f25[5]) );
  CFD2QXL \f25_reg[4]  ( .D(n208), .CP(clk), .CD(n856), .Q(f25[4]) );
  CFD2QXL \f25_reg[3]  ( .D(n206), .CP(clk), .CD(n856), .Q(f25[3]) );
  CFD2QXL \f25_reg[2]  ( .D(n204), .CP(clk), .CD(n856), .Q(f25[2]) );
  CFD2QXL \f25_reg[0]  ( .D(n202), .CP(clk), .CD(n855), .Q(f25[0]) );
  CFD2QXL \f32_reg[27]  ( .D(s32[27]), .CP(clk), .CD(n877), .Q(f32[27]) );
  CFD2QXL \f32_reg[26]  ( .D(s32[26]), .CP(clk), .CD(n877), .Q(f32[26]) );
  CFD2QXL \f32_reg[25]  ( .D(s32[25]), .CP(clk), .CD(n877), .Q(f32[25]) );
  CFD2QXL \f32_reg[24]  ( .D(s32[24]), .CP(clk), .CD(n876), .Q(f32[24]) );
  CFD2QXL \f32_reg[23]  ( .D(s32[23]), .CP(clk), .CD(n876), .Q(f32[23]) );
  CFD2QXL \f32_reg[22]  ( .D(s32[22]), .CP(clk), .CD(n876), .Q(f32[22]) );
  CFD2QXL \f32_reg[21]  ( .D(s32[21]), .CP(clk), .CD(n876), .Q(f32[21]) );
  CFD2QXL \f32_reg[20]  ( .D(s32[20]), .CP(clk), .CD(n876), .Q(f32[20]) );
  CFD2QXL \f32_reg[19]  ( .D(s32[19]), .CP(clk), .CD(n876), .Q(f32[19]) );
  CFD2QXL \f32_reg[18]  ( .D(s32[18]), .CP(clk), .CD(n875), .Q(f32[18]) );
  CFD2QXL \f32_reg[17]  ( .D(s32[17]), .CP(clk), .CD(n875), .Q(f32[17]) );
  CFD2QXL \f32_reg[16]  ( .D(s32[16]), .CP(clk), .CD(n875), .Q(f32[16]) );
  CFD2QXL \f32_reg[15]  ( .D(s32[15]), .CP(clk), .CD(n875), .Q(f32[15]) );
  CFD2QXL \f32_reg[14]  ( .D(s32[14]), .CP(clk), .CD(n875), .Q(f32[14]) );
  CFD2QXL \f32_reg[13]  ( .D(s32[13]), .CP(clk), .CD(n875), .Q(f32[13]) );
  CFD2QXL \f32_reg[12]  ( .D(s32[12]), .CP(clk), .CD(n875), .Q(f32[12]) );
  CFD2QXL \f32_reg[11]  ( .D(s32[11]), .CP(clk), .CD(n874), .Q(f32[11]) );
  CFD2QXL \f32_reg[10]  ( .D(s32[10]), .CP(clk), .CD(n874), .Q(f32[10]) );
  CFD2QXL \f32_reg[9]  ( .D(s32[9]), .CP(clk), .CD(n874), .Q(f32[9]) );
  CFD2QXL \f32_reg[8]  ( .D(s32[8]), .CP(clk), .CD(n874), .Q(f32[8]) );
  CFD2QXL \f32_reg[7]  ( .D(s32[7]), .CP(clk), .CD(n874), .Q(f32[7]) );
  CFD2QXL \f32_reg[6]  ( .D(s32[6]), .CP(clk), .CD(n874), .Q(f32[6]) );
  CFD2QXL \f32_reg[5]  ( .D(s32[5]), .CP(clk), .CD(n873), .Q(f32[5]) );
  CFD2QXL \f32_reg[4]  ( .D(s32[4]), .CP(clk), .CD(n873), .Q(f32[4]) );
  CFD2QXL \f32_reg[3]  ( .D(s32[3]), .CP(clk), .CD(n873), .Q(f32[3]) );
  CFD2QXL \f32_reg[2]  ( .D(s32[2]), .CP(clk), .CD(n873), .Q(f32[2]) );
  CFD2QXL \f32_reg[1]  ( .D(s32[1]), .CP(clk), .CD(n873), .Q(f32[1]) );
  CFD2QXL \f43_reg[27]  ( .D(s43[27]), .CP(clk), .CD(n855), .Q(f43[27]) );
  CFD2QXL \f43_reg[26]  ( .D(s43[26]), .CP(clk), .CD(n855), .Q(f43[26]) );
  CFD2QXL \f43_reg[25]  ( .D(s43[25]), .CP(clk), .CD(n854), .Q(f43[25]) );
  CFD2QXL \f43_reg[24]  ( .D(s43[24]), .CP(clk), .CD(n854), .Q(f43[24]) );
  CFD2QXL \f43_reg[23]  ( .D(s43[23]), .CP(clk), .CD(n854), .Q(f43[23]) );
  CFD2QXL \f43_reg[22]  ( .D(s43[22]), .CP(clk), .CD(n854), .Q(f43[22]) );
  CFD2QXL \f43_reg[21]  ( .D(s43[21]), .CP(clk), .CD(n854), .Q(f43[21]) );
  CFD2QXL \f43_reg[20]  ( .D(s43[20]), .CP(clk), .CD(n854), .Q(f43[20]) );
  CFD2QXL \f43_reg[19]  ( .D(s43[19]), .CP(clk), .CD(n853), .Q(f43[19]) );
  CFD2QXL \f43_reg[18]  ( .D(s43[18]), .CP(clk), .CD(n853), .Q(f43[18]) );
  CFD2QXL \f43_reg[17]  ( .D(s43[17]), .CP(clk), .CD(n853), .Q(f43[17]) );
  CFD2QXL \f43_reg[16]  ( .D(s43[16]), .CP(clk), .CD(n853), .Q(f43[16]) );
  CFD2QXL \f43_reg[15]  ( .D(s43[15]), .CP(clk), .CD(n853), .Q(f43[15]) );
  CFD2QXL \f43_reg[14]  ( .D(s43[14]), .CP(clk), .CD(n853), .Q(f43[14]) );
  CFD2QXL \f43_reg[13]  ( .D(s43[13]), .CP(clk), .CD(n853), .Q(f43[13]) );
  CFD2QXL \f43_reg[12]  ( .D(s43[12]), .CP(clk), .CD(n852), .Q(f43[12]) );
  CFD2QXL \f43_reg[11]  ( .D(s43[11]), .CP(clk), .CD(n852), .Q(f43[11]) );
  CFD2QXL \f43_reg[10]  ( .D(s43[10]), .CP(clk), .CD(n852), .Q(f43[10]) );
  CFD2QXL \f43_reg[9]  ( .D(s43[9]), .CP(clk), .CD(n852), .Q(f43[9]) );
  CFD2QXL \f43_reg[8]  ( .D(s43[8]), .CP(clk), .CD(n852), .Q(f43[8]) );
  CFD2QXL \f43_reg[7]  ( .D(s43[7]), .CP(clk), .CD(n852), .Q(f43[7]) );
  CFD2QXL \f43_reg[6]  ( .D(s43[6]), .CP(clk), .CD(n851), .Q(f43[6]) );
  CFD2QXL \f43_reg[5]  ( .D(s43[5]), .CP(clk), .CD(n851), .Q(f43[5]) );
  CFD2QXL \f43_reg[4]  ( .D(s43[4]), .CP(clk), .CD(n851), .Q(f43[4]) );
  CFD2QXL \f43_reg[3]  ( .D(s43[3]), .CP(clk), .CD(n851), .Q(f43[3]) );
  CFD2QXL \f43_reg[2]  ( .D(s43[2]), .CP(clk), .CD(n851), .Q(f43[2]) );
  CFD2QXL \res_d_reg[1]  ( .D(res_temp[1]), .CP(clk), .CD(n850), .Q(res_d[1])
         );
  CFD2QXL \res_d_reg[2]  ( .D(res_temp[2]), .CP(clk), .CD(n850), .Q(res_d[2])
         );
  CFD2QXL \res_d_reg[3]  ( .D(res_temp[3]), .CP(clk), .CD(n850), .Q(res_d[3])
         );
  CFD2QXL \res_d_reg[4]  ( .D(res_temp[4]), .CP(clk), .CD(n850), .Q(res_d[4])
         );
  CFD2QXL \res_d_reg[5]  ( .D(res_temp[5]), .CP(clk), .CD(n850), .Q(res_d[5])
         );
  CFD2QXL \res_d_reg[6]  ( .D(res_temp[6]), .CP(clk), .CD(n849), .Q(res_d[6])
         );
  CFD2QXL \res_d_reg[7]  ( .D(res_temp[7]), .CP(clk), .CD(n849), .Q(res_d[7])
         );
  CFD2QXL \res_d_reg[8]  ( .D(res_temp[8]), .CP(clk), .CD(n849), .Q(res_d[8])
         );
  CFD2QXL \res_d_reg[9]  ( .D(res_temp[9]), .CP(clk), .CD(n849), .Q(res_d[9])
         );
  CFD2QXL \res_d_reg[10]  ( .D(res_temp[10]), .CP(clk), .CD(n849), .Q(
        res_d[10]) );
  CFD2QXL \res_d_reg[11]  ( .D(res_temp[11]), .CP(clk), .CD(n849), .Q(
        res_d[11]) );
  CFD2QXL \res_d_reg[12]  ( .D(res_temp[12]), .CP(clk), .CD(n849), .Q(
        res_d[12]) );
  CFD2QXL \res_d_reg[13]  ( .D(res_temp[13]), .CP(clk), .CD(n848), .Q(
        res_d[13]) );
  CFD2QXL \res_d_reg[14]  ( .D(res_temp[14]), .CP(clk), .CD(n848), .Q(
        res_d[14]) );
  CFD2QXL \res_d_reg[15]  ( .D(res_temp[15]), .CP(clk), .CD(n848), .Q(
        res_d[15]) );
  CFD2QXL \res_d_reg[16]  ( .D(res_temp[16]), .CP(clk), .CD(n848), .Q(
        res_d[16]) );
  CFD2QXL \res_d_reg[17]  ( .D(res_temp[17]), .CP(clk), .CD(n848), .Q(
        res_d[17]) );
  CFD2QXL \res_d_reg[18]  ( .D(res_temp[18]), .CP(clk), .CD(n848), .Q(
        res_d[18]) );
  CFD2QXL \res_d_reg[19]  ( .D(res_temp[19]), .CP(clk), .CD(n847), .Q(
        res_d[19]) );
  CFD2QXL \res_d_reg[20]  ( .D(res_temp[20]), .CP(clk), .CD(n847), .Q(
        res_d[20]) );
  CFD2QXL \res_d_reg[21]  ( .D(res_temp[21]), .CP(clk), .CD(n847), .Q(
        res_d[21]) );
  CFD2QXL \res_d_reg[22]  ( .D(res_temp[22]), .CP(clk), .CD(n847), .Q(
        res_d[22]) );
  CFD2QXL \res_d_reg[23]  ( .D(res_temp[23]), .CP(clk), .CD(n847), .Q(
        res_d[23]) );
  CFD2QXL \res_d_reg[24]  ( .D(res_temp[24]), .CP(clk), .CD(n847), .Q(
        res_d[24]) );
  CFD2QXL \res_d_reg[25]  ( .D(res_temp[25]), .CP(clk), .CD(n847), .Q(
        res_d[25]) );
  CFD2QXL \res_d_reg[26]  ( .D(res_temp[26]), .CP(clk), .CD(n846), .Q(
        res_d[26]) );
  CFD2QXL \res_d_reg[27]  ( .D(res_temp[27]), .CP(clk), .CD(n846), .Q(
        res_d[27]) );
  CFD2QXL pushOut_reg ( .D(n200), .CP(clk), .CD(n925), .Q(pushZ) );
  CFD2QXL \res_reg[0]  ( .D(n198), .CP(clk), .CD(n850), .Q(Z[0]) );
  CFD2QXL \res_reg[1]  ( .D(n196), .CP(clk), .CD(n850), .Q(Z[1]) );
  CFD2QXL \res_reg[2]  ( .D(n194), .CP(clk), .CD(n850), .Q(Z[2]) );
  CFD2QXL \res_reg[3]  ( .D(n192), .CP(clk), .CD(n850), .Q(Z[3]) );
  CFD2QXL \res_reg[4]  ( .D(n190), .CP(clk), .CD(n850), .Q(Z[4]) );
  CFD2QXL \res_reg[5]  ( .D(n188), .CP(clk), .CD(n850), .Q(Z[5]) );
  CFD2QXL \res_reg[6]  ( .D(n186), .CP(clk), .CD(n849), .Q(Z[6]) );
  CFD2QXL \res_reg[7]  ( .D(n184), .CP(clk), .CD(n849), .Q(Z[7]) );
  CFD2QXL \res_reg[8]  ( .D(n182), .CP(clk), .CD(n849), .Q(Z[8]) );
  CFD2QXL \res_reg[9]  ( .D(n180), .CP(clk), .CD(n849), .Q(Z[9]) );
  CFD2QXL \res_reg[10]  ( .D(n178), .CP(clk), .CD(n849), .Q(Z[10]) );
  CFD2QXL \res_reg[11]  ( .D(n176), .CP(clk), .CD(n849), .Q(Z[11]) );
  CFD2QXL \res_reg[12]  ( .D(n174), .CP(clk), .CD(n848), .Q(Z[12]) );
  CFD2QXL \res_reg[13]  ( .D(n172), .CP(clk), .CD(n848), .Q(Z[13]) );
  CFD2QXL \res_reg[14]  ( .D(n170), .CP(clk), .CD(n848), .Q(Z[14]) );
  CFD2QXL \res_reg[15]  ( .D(n168), .CP(clk), .CD(n848), .Q(Z[15]) );
  CFD2QXL \res_reg[16]  ( .D(n166), .CP(clk), .CD(n848), .Q(Z[16]) );
  CFD2QXL \res_reg[17]  ( .D(n164), .CP(clk), .CD(n848), .Q(Z[17]) );
  CFD2QXL \res_reg[18]  ( .D(n162), .CP(clk), .CD(n848), .Q(Z[18]) );
  CFD2QXL \res_reg[19]  ( .D(n160), .CP(clk), .CD(n847), .Q(Z[19]) );
  CFD2QXL \res_reg[20]  ( .D(n158), .CP(clk), .CD(n847), .Q(Z[20]) );
  CFD2QXL \res_reg[21]  ( .D(n156), .CP(clk), .CD(n847), .Q(Z[21]) );
  CFD2QXL \res_reg[22]  ( .D(n154), .CP(clk), .CD(n847), .Q(Z[22]) );
  CFD2QXL \res_reg[23]  ( .D(n152), .CP(clk), .CD(n847), .Q(Z[23]) );
  CFD2QXL \res_reg[24]  ( .D(n150), .CP(clk), .CD(n847), .Q(Z[24]) );
  CFD2QXL \res_reg[25]  ( .D(n148), .CP(clk), .CD(n846), .Q(Z[25]) );
  CFD2QXL \res_reg[26]  ( .D(n146), .CP(clk), .CD(n846), .Q(Z[26]) );
  CFD2QXL \res_reg[27]  ( .D(n144), .CP(clk), .CD(n846), .Q(Z[27]) );
  CFD2QXL \res_reg[28]  ( .D(n142), .CP(clk), .CD(n846), .Q(Z[28]) );
  CFD2QXL \res_reg[29]  ( .D(n140), .CP(clk), .CD(n846), .Q(Z[29]) );
  CFD2QXL \res_reg[30]  ( .D(n138), .CP(clk), .CD(n846), .Q(Z[30]) );
  CFD2QXL \res_reg[31]  ( .D(n136), .CP(clk), .CD(n846), .Q(Z[31]) );
  CFD2QXL \f23_reg[25]  ( .D(s23[25]), .CP(clk), .CD(n914), .Q(f23[25]) );
  CFD2QXL \f31_reg[23]  ( .D(s31[23]), .CP(clk), .CD(n909), .Q(f31[23]) );
  CFD2QXL \f21_reg[13]  ( .D(n135), .CP(clk), .CD(n911), .Q(f21[13]) );
  CFD2QXL \f21_reg[10]  ( .D(n133), .CP(clk), .CD(n910), .Q(f21[10]) );
  CFD2QXL \f21_reg[8]  ( .D(n131), .CP(clk), .CD(n910), .Q(f21[8]) );
  CFD2QXL \f21_reg[6]  ( .D(n129), .CP(clk), .CD(n910), .Q(f21[6]) );
  CFD2QXL \f14_reg[0]  ( .D(s14[0]), .CP(clk), .CD(n892), .Q(f14[0]) );
  CFD2QXL \f13_reg[29]  ( .D(n572), .CP(clk), .CD(n901), .Q(f13[29]) );
  CFD2QX1 \f11_reg[8]  ( .D(n826), .CP(clk), .CD(n915), .Q(f11[8]) );
  CFD2QX1 \f13_reg[8]  ( .D(n122), .CP(clk), .CD(n897), .Q(f13[8]) );
  CFD2QX1 \f02_reg[20]  ( .D(n824), .CP(clk), .CD(n899), .Q(f02[20]) );
  CFD2QX1 \f02_reg[24]  ( .D(n823), .CP(clk), .CD(n900), .Q(f02[24]) );
  CFD2QX1 \f01_reg[18]  ( .D(n822), .CP(clk), .CD(n922), .Q(f01[18]) );
  CFD2QX1 \f31_reg[0]  ( .D(s31[0]), .CP(clk), .CD(n907), .Q(f31[0]) );
  CFD2QXL \f14_reg[12]  ( .D(s14[12]), .CP(clk), .CD(n893), .Q(f14[12]) );
  CFD2QXL \f30_reg[14]  ( .D(n662), .CP(clk), .CD(n906), .Q(f30[14]) );
  CFD2QXL \f30_reg[13]  ( .D(n661), .CP(clk), .CD(n906), .Q(f30[13]) );
  CFD2QXL \f30_reg[1]  ( .D(n659), .CP(clk), .CD(n905), .Q(f30[1]) );
  CFD2QX1 \f17_reg[5]  ( .D(s17[5]), .CP(clk), .CD(n880), .Q(f17[5]) );
  CFD2QXL \f30_reg[19]  ( .D(n821), .CP(clk), .CD(n906), .Q(f30[19]) );
  CFD2QX1 \f31_reg[1]  ( .D(s31[1]), .CP(clk), .CD(n907), .Q(f31[1]) );
  CFD2QX1 \f03_reg[24]  ( .D(n723), .CP(clk), .CD(n889), .Q(f03[24]) );
  CFD2QXL \f30_reg[20]  ( .D(f21[20]), .CP(clk), .CD(n906), .Q(f30[20]) );
  CFD2QXL \f11_reg[29]  ( .D(n664), .CP(clk), .CD(n917), .Q(f11[29]) );
  CFD2QXL \f30_reg[0]  ( .D(n814), .CP(clk), .CD(n905), .Q(f30[0]) );
  CFD2QX1 \f11_reg[0]  ( .D(n696), .CP(clk), .CD(n914), .Q(f11[0]) );
  CFD2QX1 \f11_reg[4]  ( .D(n447), .CP(clk), .CD(n915), .Q(f11[4]) );
  CFD2QX1 \f12_reg[11]  ( .D(s12[11]), .CP(clk), .CD(n918), .Q(f12[11]) );
  CFD2QXL \f14_reg[2]  ( .D(s14[2]), .CP(clk), .CD(n892), .Q(f14[2]) );
  CFD2QXL \f14_reg[14]  ( .D(s14[14]), .CP(clk), .CD(n893), .Q(f14[14]) );
  CFD2QXL \f14_reg[13]  ( .D(s14[13]), .CP(clk), .CD(n893), .Q(f14[13]) );
  CFD2QXL \f14_reg[10]  ( .D(s14[10]), .CP(clk), .CD(n893), .Q(f14[10]) );
  CFD2QXL \f14_reg[11]  ( .D(s14[11]), .CP(clk), .CD(n893), .Q(f14[11]) );
  CFD2QXL \f14_reg[8]  ( .D(s14[8]), .CP(clk), .CD(n893), .Q(f14[8]) );
  CFD2QXL \f14_reg[6]  ( .D(s14[6]), .CP(clk), .CD(n893), .Q(f14[6]) );
  CFD2QXL \f14_reg[4]  ( .D(s14[4]), .CP(clk), .CD(n893), .Q(f14[4]) );
  CFD2QXL \f14_reg[3]  ( .D(s14[3]), .CP(clk), .CD(n893), .Q(f14[3]) );
  CFD2QXL \f17_reg[8]  ( .D(s17[8]), .CP(clk), .CD(n881), .Q(f17[8]) );
  CFD2QXL \f17_reg[13]  ( .D(s17[13]), .CP(clk), .CD(n881), .Q(f17[13]) );
  CFD2QXL \f17_reg[11]  ( .D(s17[11]), .CP(clk), .CD(n881), .Q(f17[11]) );
  CFD2QXL \f17_reg[9]  ( .D(s17[9]), .CP(clk), .CD(n881), .Q(f17[9]) );
  CFD2QXL \f17_reg[7]  ( .D(s17[7]), .CP(clk), .CD(n881), .Q(f17[7]) );
  CFD2QXL \f17_reg[6]  ( .D(s17[6]), .CP(clk), .CD(n880), .Q(f17[6]) );
  CFD2QXL \f17_reg[12]  ( .D(s17[12]), .CP(clk), .CD(n881), .Q(f17[12]) );
  CFD2QXL \f17_reg[10]  ( .D(s17[10]), .CP(clk), .CD(n881), .Q(f17[10]) );
  CFD2QXL \f23_reg[16]  ( .D(s23[16]), .CP(clk), .CD(n913), .Q(f23[16]) );
  CFD2QXL \f23_reg[0]  ( .D(s23[0]), .CP(clk), .CD(n912), .Q(f23[0]) );
  CFD2QXL \f31_reg[12]  ( .D(s31[12]), .CP(clk), .CD(n908), .Q(f31[12]) );
  CFD2QXL \f14_reg[18]  ( .D(s14[18]), .CP(clk), .CD(n894), .Q(f14[18]) );
  CFD2QXL \f17_reg[16]  ( .D(s17[16]), .CP(clk), .CD(n881), .Q(f17[16]) );
  CFD2QXL \f03_reg[25]  ( .D(n670), .CP(clk), .CD(n889), .Q(f03[25]) );
  CFD2QX1 \f23_reg[3]  ( .D(s23[3]), .CP(clk), .CD(n912), .Q(f23[3]) );
  CFD2QX2 \f11_reg[7]  ( .D(n668), .CP(clk), .CD(n915), .Q(f11[7]) );
  CFD2QX1 \f23_reg[12]  ( .D(s23[12]), .CP(clk), .CD(n913), .Q(f23[12]) );
  CFD2QX1 \f12_reg[15]  ( .D(s12[15]), .CP(clk), .CD(n918), .Q(f12[15]) );
  CFD2QX1 \f11_reg[5]  ( .D(n650), .CP(clk), .CD(n915), .Q(f11[5]) );
  CFD2QX2 \f02_reg[10]  ( .D(n648), .CP(clk), .CD(n897), .Q(f02[10]) );
  CFD2QX1 \f01_reg[14]  ( .D(n647), .CP(clk), .CD(n922), .Q(f01[14]) );
  CFD2QX2 \f12_reg[13]  ( .D(s12[13]), .CP(clk), .CD(n918), .Q(f12[13]) );
  CFD2QX1 \f12_reg[17]  ( .D(s12[17]), .CP(clk), .CD(n918), .Q(f12[17]) );
  CFD2QX1 \f12_reg[9]  ( .D(s12[9]), .CP(clk), .CD(n918), .Q(f12[9]) );
  CFD2QX1 \f03_reg[23]  ( .D(n641), .CP(clk), .CD(n888), .Q(f03[23]) );
  CFD2QX1 \f31_reg[2]  ( .D(s31[2]), .CP(clk), .CD(n907), .Q(f31[2]) );
  CFD2QX1 \f13_reg[28]  ( .D(n640), .CP(clk), .CD(n901), .Q(f13[28]) );
  CFD2QX1 \f17_reg[15]  ( .D(s17[15]), .CP(clk), .CD(n881), .Q(f17[15]) );
  CFD2QX1 \f02_reg[29]  ( .D(n639), .CP(clk), .CD(n902), .Q(f02[29]) );
  CFD2QX1 \f01_reg[29]  ( .D(n638), .CP(clk), .CD(n924), .Q(f01[29]) );
  CFD2QX1 \f01_reg[20]  ( .D(n637), .CP(clk), .CD(n922), .Q(f01[20]) );
  CFD2QX1 \f02_reg[9]  ( .D(n636), .CP(clk), .CD(n897), .Q(f02[9]) );
  CFD2QX1 \f02_reg[17]  ( .D(n635), .CP(clk), .CD(n899), .Q(f02[17]) );
  CFD2QX1 \f02_reg[6]  ( .D(n628), .CP(clk), .CD(n896), .Q(f02[6]) );
  CFD2QX1 \f13_reg[10]  ( .D(n627), .CP(clk), .CD(n897), .Q(f13[10]) );
  CFD2QX1 \f02_reg[26]  ( .D(n626), .CP(clk), .CD(n901), .Q(f02[26]) );
  CFD2QX1 \f01_reg[15]  ( .D(n624), .CP(clk), .CD(n922), .Q(f01[15]) );
  CFD2QX1 \f21_reg[16]  ( .D(n614), .CP(clk), .CD(n911), .Q(f21[16]) );
  CFD2QX1 \f13_reg[9]  ( .D(n612), .CP(clk), .CD(n897), .Q(f13[9]) );
  CFD2QX1 \f01_reg[16]  ( .D(n611), .CP(clk), .CD(n922), .Q(f01[16]) );
  CFD2QX2 \f11_reg[16]  ( .D(n606), .CP(clk), .CD(n916), .Q(f11[16]) );
  CFD2QX1 \f02_reg[19]  ( .D(n607), .CP(clk), .CD(n899), .Q(f02[19]) );
  CFD2QX1 \f13_reg[19]  ( .D(n608), .CP(clk), .CD(n899), .Q(f13[19]) );
  CFD2QX1 \f11_reg[26]  ( .D(n604), .CP(clk), .CD(n916), .Q(f11[26]) );
  CFD2QX1 \f31_reg[21]  ( .D(s31[21]), .CP(clk), .CD(n909), .Q(f31[21]) );
  CFD2QX1 \f23_reg[11]  ( .D(s23[11]), .CP(clk), .CD(n913), .Q(f23[11]) );
  CFD2QX1 \f11_reg[3]  ( .D(n691), .CP(clk), .CD(n915), .Q(f11[3]) );
  CFD2QX1 \f11_reg[25]  ( .D(n655), .CP(clk), .CD(n916), .Q(f11[25]) );
  CFD2QX1 \f01_reg[21]  ( .D(n654), .CP(clk), .CD(n923), .Q(f01[21]) );
  CFD2QX1 \f11_reg[21]  ( .D(n651), .CP(clk), .CD(n916), .Q(f11[21]) );
  CFD2QX1 \f23_reg[19]  ( .D(s23[19]), .CP(clk), .CD(n913), .Q(f23[19]) );
  CFD2QX1 \f31_reg[14]  ( .D(s31[14]), .CP(clk), .CD(n908), .Q(f31[14]) );
  CFD2QX1 \f01_reg[22]  ( .D(n629), .CP(clk), .CD(n923), .Q(f01[22]) );
  CFD2QX1 \f01_reg[26]  ( .D(n617), .CP(clk), .CD(n923), .Q(f01[26]) );
  CFD2QX1 \f13_reg[0]  ( .D(n693), .CP(clk), .CD(n895), .Q(f13[0]) );
  CFD2QX1 \f13_reg[20]  ( .D(n710), .CP(clk), .CD(n899), .Q(f13[20]) );
  CFD2QX1 \f01_reg[24]  ( .D(n681), .CP(clk), .CD(n923), .Q(f01[24]) );
  CFD2QX1 \f23_reg[20]  ( .D(s23[20]), .CP(clk), .CD(n914), .Q(f23[20]) );
  CFD2QX1 \f11_reg[6]  ( .D(n622), .CP(clk), .CD(n915), .Q(f11[6]) );
  CFD2QX1 \f31_reg[19]  ( .D(s31[19]), .CP(clk), .CD(n909), .Q(f31[19]) );
  CFD2QX1 \f30_reg[16]  ( .D(n618), .CP(clk), .CD(n906), .Q(f30[16]) );
  CFD2QX1 \f31_reg[11]  ( .D(s31[11]), .CP(clk), .CD(n908), .Q(f31[11]) );
  CFD2QX1 \f17_reg[0]  ( .D(s17[0]), .CP(clk), .CD(n880), .Q(f17[0]) );
  CFD2QX1 \f30_reg[17]  ( .D(n687), .CP(clk), .CD(n906), .Q(f30[17]) );
  CFD2QX1 \f23_reg[6]  ( .D(s23[6]), .CP(clk), .CD(n912), .Q(f23[6]) );
  CFD2QX1 \f23_reg[17]  ( .D(s23[17]), .CP(clk), .CD(n913), .Q(f23[17]) );
  CFD2QX1 \f12_reg[23]  ( .D(s12[23]), .CP(clk), .CD(n919), .Q(f12[23]) );
  CFD2QX1 \f17_reg[18]  ( .D(s17[18]), .CP(clk), .CD(n881), .Q(f17[18]) );
  CFD2QX1 \f31_reg[15]  ( .D(s31[15]), .CP(clk), .CD(n908), .Q(f31[15]) );
  CFD2QX1 \f31_reg[16]  ( .D(s31[16]), .CP(clk), .CD(n908), .Q(f31[16]) );
  CFD2QX1 \f31_reg[3]  ( .D(s31[3]), .CP(clk), .CD(n907), .Q(f31[3]) );
  CFD2QX1 \f14_reg[20]  ( .D(s14[20]), .CP(clk), .CD(n894), .Q(f14[20]) );
  CFD2QX1 \f23_reg[18]  ( .D(s23[18]), .CP(clk), .CD(n913), .Q(f23[18]) );
  CFD2QX1 \f31_reg[10]  ( .D(s31[10]), .CP(clk), .CD(n908), .Q(f31[10]) );
  CFD2QX1 \f17_reg[3]  ( .D(s17[3]), .CP(clk), .CD(n880), .Q(f17[3]) );
  CFD2QX1 \f31_reg[4]  ( .D(s31[4]), .CP(clk), .CD(n907), .Q(f31[4]) );
  CFD2QX1 \f23_reg[4]  ( .D(s23[4]), .CP(clk), .CD(n912), .Q(f23[4]) );
  CFD2QX1 \f01_reg[5]  ( .D(n574), .CP(clk), .CD(n920), .Q(f01[5]) );
  CFD2QX2 \f11_reg[17]  ( .D(n678), .CP(clk), .CD(n916), .Q(f11[17]) );
  CFD2QX1 \f01_reg[17]  ( .D(n682), .CP(clk), .CD(n922), .Q(f01[17]) );
  CFD2QX1 \f02_reg[22]  ( .D(n674), .CP(clk), .CD(n900), .Q(f02[22]) );
  CFD2QX1 \f14_reg[19]  ( .D(s14[19]), .CP(clk), .CD(n894), .Q(f14[19]) );
  CFD2QX2 \f11_reg[15]  ( .D(n833), .CP(clk), .CD(n916), .Q(f11[15]) );
  CFD2QX2 \f11_reg[22]  ( .D(n675), .CP(clk), .CD(n916), .Q(f11[22]) );
  CFD2QX1 \f17_reg[19]  ( .D(s17[19]), .CP(clk), .CD(n881), .Q(f17[19]) );
  CFD2QX1 \f21_reg[0]  ( .D(n564), .CP(clk), .CD(n910), .Q(f21[0]) );
  CFD2QX1 \f23_reg[2]  ( .D(s23[2]), .CP(clk), .CD(n912), .Q(f23[2]) );
  CFD2QX1 \f17_reg[4]  ( .D(s17[4]), .CP(clk), .CD(n880), .Q(f17[4]) );
  CFD2QX1 \f11_reg[9]  ( .D(n790), .CP(clk), .CD(n915), .Q(f11[9]) );
  CFD2QXL \f21_reg[1]  ( .D(n688), .CP(clk), .CD(n910), .Q(f21[1]) );
  CFD2QX1 \f23_reg[1]  ( .D(s23[1]), .CP(clk), .CD(n912), .Q(f23[1]) );
  CFD2QX1 \f23_reg[21]  ( .D(s23[21]), .CP(clk), .CD(n914), .Q(f23[21]) );
  CFD2QX1 \f31_reg[25]  ( .D(s31[25]), .CP(clk), .CD(n909), .Q(f31[25]) );
  CFD2QX1 \f30_reg[18]  ( .D(n120), .CP(clk), .CD(n906), .Q(f30[18]) );
  CFD2QX1 \f17_reg[17]  ( .D(s17[17]), .CP(clk), .CD(n881), .Q(f17[17]) );
  CFD2QX1 \f03_reg[26]  ( .D(n667), .CP(clk), .CD(n889), .Q(f03[26]) );
  CFD2QX1 \f31_reg[13]  ( .D(s31[13]), .CP(clk), .CD(n908), .Q(f31[13]) );
  CFD2QX2 \f11_reg[23]  ( .D(n642), .CP(clk), .CD(n916), .Q(f11[23]) );
  CFD2QX1 \f11_reg[19]  ( .D(n665), .CP(clk), .CD(n916), .Q(f11[19]) );
  CFD2QX1 \f12_reg[5]  ( .D(s12[5]), .CP(clk), .CD(n917), .Q(f12[5]) );
  CFD2QX1 \f12_reg[0]  ( .D(s12[0]), .CP(clk), .CD(n917), .Q(f12[0]) );
  CFD2QX1 \f17_reg[2]  ( .D(s17[2]), .CP(clk), .CD(n880), .Q(f17[2]) );
  CFD2QX1 \f01_reg[27]  ( .D(n819), .CP(clk), .CD(n924), .Q(f01[27]) );
  CFD2QX1 \f31_reg[29]  ( .D(s31[29]), .CP(clk), .CD(n909), .Q(f31[29]) );
  CFD2QX1 \f03_reg[5]  ( .D(n580), .CP(clk), .CD(n886), .Q(f03[5]) );
  CFD2QX1 \f23_reg[7]  ( .D(s23[7]), .CP(clk), .CD(n913), .Q(f23[7]) );
  CFD2QX1 \f01_reg[7]  ( .D(n804), .CP(clk), .CD(n920), .Q(f01[7]) );
  CFD2QX1 \f03_reg[3]  ( .D(n738), .CP(clk), .CD(n885), .Q(f03[3]) );
  CFD2QX1 \f02_reg[13]  ( .D(n780), .CP(clk), .CD(n898), .Q(f02[13]) );
  CFD2QX1 \f03_reg[4]  ( .D(n577), .CP(clk), .CD(n886), .Q(f03[4]) );
  CFD2QX1 \f03_reg[2]  ( .D(n736), .CP(clk), .CD(n885), .Q(f03[2]) );
  CFD2QX1 \f01_reg[3]  ( .D(n800), .CP(clk), .CD(n920), .Q(f01[3]) );
  CFD2QX1 \f03_reg[1]  ( .D(n734), .CP(clk), .CD(n885), .Q(f03[1]) );
  CFD2QX2 \f03_reg[9]  ( .D(n598), .CP(clk), .CD(n886), .Q(f03[9]) );
  CFD2QX1 \f01_reg[1]  ( .D(n796), .CP(clk), .CD(n920), .Q(f01[1]) );
  CFD2QX1 \f01_reg[6]  ( .D(n645), .CP(clk), .CD(n920), .Q(f01[6]) );
  CFD2QX1 \f01_reg[11]  ( .D(n812), .CP(clk), .CD(n921), .Q(f01[11]) );
  CFD2QX1 \f02_reg[1]  ( .D(n762), .CP(clk), .CD(n895), .Q(f02[1]) );
  CFD2QX1 \f12_reg[7]  ( .D(s12[7]), .CP(clk), .CD(n917), .Q(f12[7]) );
  CFD2QX1 \f12_reg[2]  ( .D(s12[2]), .CP(clk), .CD(n917), .Q(f12[2]) );
  CFD2QX1 \f01_reg[10]  ( .D(n810), .CP(clk), .CD(n921), .Q(f01[10]) );
  CFD2QX1 \f01_reg[9]  ( .D(n808), .CP(clk), .CD(n921), .Q(f01[9]) );
  CFD2QX1 \f01_reg[8]  ( .D(n806), .CP(clk), .CD(n921), .Q(f01[8]) );
  CFD2QX1 \f01_reg[4]  ( .D(n802), .CP(clk), .CD(n920), .Q(f01[4]) );
  CFD2QX1 \f01_reg[2]  ( .D(n798), .CP(clk), .CD(n920), .Q(f01[2]) );
  CFD2QX1 \f02_reg[18]  ( .D(n788), .CP(clk), .CD(n899), .Q(f02[18]) );
  CFD2QX1 \f02_reg[16]  ( .D(n786), .CP(clk), .CD(n899), .Q(f02[16]) );
  CFD2QX1 \f02_reg[14]  ( .D(n782), .CP(clk), .CD(n898), .Q(f02[14]) );
  CFD2QX1 \f02_reg[12]  ( .D(n778), .CP(clk), .CD(n898), .Q(f02[12]) );
  CFD2QX1 \f02_reg[4]  ( .D(n768), .CP(clk), .CD(n896), .Q(f02[4]) );
  CFD2QX1 \f02_reg[2]  ( .D(n764), .CP(clk), .CD(n895), .Q(f02[2]) );
  CFD2QX1 \f02_reg[0]  ( .D(n760), .CP(clk), .CD(n895), .Q(f02[0]) );
  CFD2QX1 \f03_reg[22]  ( .D(n758), .CP(clk), .CD(n888), .Q(f03[22]) );
  CFD2QX1 \f03_reg[21]  ( .D(n756), .CP(clk), .CD(n888), .Q(f03[21]) );
  CFD2QX1 \f03_reg[20]  ( .D(n754), .CP(clk), .CD(n888), .Q(f03[20]) );
  CFD2QX1 \f03_reg[19]  ( .D(n752), .CP(clk), .CD(n888), .Q(f03[19]) );
  CFD2QX1 \f11_reg[27]  ( .D(n731), .CP(clk), .CD(n917), .Q(f11[27]) );
  CFD2QX1 \f11_reg[24]  ( .D(n729), .CP(clk), .CD(n916), .Q(f11[24]) );
  CFD2QX1 \f11_reg[18]  ( .D(n727), .CP(clk), .CD(n916), .Q(f11[18]) );
  CFD2QX1 \f11_reg[10]  ( .D(n726), .CP(clk), .CD(n915), .Q(f11[10]) );
  CFD2QX1 \f12_reg[28]  ( .D(s12[28]), .CP(clk), .CD(n919), .Q(f12[28]) );
  CFD2QX1 \f12_reg[8]  ( .D(s12[8]), .CP(clk), .CD(n918), .Q(f12[8]) );
  CFD2QX1 \f12_reg[6]  ( .D(s12[6]), .CP(clk), .CD(n917), .Q(f12[6]) );
  CFD2QX1 \f13_reg[24]  ( .D(n717), .CP(clk), .CD(n900), .Q(f13[24]) );
  CFD2QX1 \f13_reg[22]  ( .D(n712), .CP(clk), .CD(n900), .Q(f13[22]) );
  CFD2QX1 \f13_reg[2]  ( .D(n702), .CP(clk), .CD(n895), .Q(f13[2]) );
  CFD2QX1 \f23_reg[8]  ( .D(s23[8]), .CP(clk), .CD(n913), .Q(f23[8]) );
  CFD2QX2 \f03_reg[15]  ( .D(n594), .CP(clk), .CD(n887), .Q(f03[15]) );
  CFD2QX1 \f31_reg[6]  ( .D(s31[6]), .CP(clk), .CD(n908), .Q(f31[6]) );
  CFD2QX1 \f01_reg[12]  ( .D(n632), .CP(clk), .CD(n921), .Q(f01[12]) );
  CFD2QX2 \f03_reg[16]  ( .D(n615), .CP(clk), .CD(n887), .Q(f03[16]) );
  CFD2QX1 \f13_reg[4]  ( .D(n694), .CP(clk), .CD(n896), .Q(f13[4]) );
  CFD2QX1 \f17_reg[14]  ( .D(s17[14]), .CP(clk), .CD(n881), .Q(f17[14]) );
  CFD2QX1 \f12_reg[26]  ( .D(s12[26]), .CP(clk), .CD(n919), .Q(f12[26]) );
  CFD2QX1 \f12_reg[16]  ( .D(s12[16]), .CP(clk), .CD(n918), .Q(f12[16]) );
  CFD2QX1 \f12_reg[22]  ( .D(s12[22]), .CP(clk), .CD(n919), .Q(f12[22]) );
  CFD2QX1 \f13_reg[6]  ( .D(n634), .CP(clk), .CD(n896), .Q(f13[6]) );
  CFD2QX1 \f13_reg[26]  ( .D(n119), .CP(clk), .CD(n901), .Q(f13[26]) );
  CFD2QX1 \f02_reg[23]  ( .D(n620), .CP(clk), .CD(n900), .Q(f02[23]) );
  CFD2QX1 \f02_reg[25]  ( .D(n602), .CP(clk), .CD(n901), .Q(f02[25]) );
  CFD2QX1 \f01_reg[25]  ( .D(n657), .CP(clk), .CD(n923), .Q(f01[25]) );
  CFD2QX2 \f11_reg[14]  ( .D(n630), .CP(clk), .CD(n916), .Q(f11[14]) );
  CFD2QX1 \f23_reg[24]  ( .D(s23[24]), .CP(clk), .CD(n914), .Q(f23[24]) );
  CFD2QXL \f23_reg[10]  ( .D(s23[10]), .CP(clk), .CD(n913), .Q(f23[10]) );
  CFD2QX1 \f23_reg[22]  ( .D(s23[22]), .CP(clk), .CD(n914), .Q(f23[22]) );
  CFD2QXL \f31_reg[20]  ( .D(s31[20]), .CP(clk), .CD(n909), .Q(f31[20]) );
  CFD2QXL \f31_reg[18]  ( .D(s31[18]), .CP(clk), .CD(n908), .Q(f31[18]) );
  CFD2QX1 \f31_reg[17]  ( .D(s31[17]), .CP(clk), .CD(n908), .Q(f31[17]) );
  CFD2QX2 \f03_reg[7]  ( .D(n817), .CP(clk), .CD(n886), .Q(f03[7]) );
  CFD2QX1 \f31_reg[22]  ( .D(s31[22]), .CP(clk), .CD(n909), .Q(f31[22]) );
  CFD2QX1 \f31_reg[24]  ( .D(s31[24]), .CP(clk), .CD(n909), .Q(f31[24]) );
  CFD2QXL \f14_reg[16]  ( .D(s14[16]), .CP(clk), .CD(n894), .Q(f14[16]) );
  CFD2QX1 \f01_reg[23]  ( .D(n685), .CP(clk), .CD(n923), .Q(f01[23]) );
  CFD2QXL \f31_reg[8]  ( .D(s31[8]), .CP(clk), .CD(n908), .Q(f31[8]) );
  CFD2QX1 \f11_reg[1]  ( .D(n683), .CP(clk), .CD(n915), .Q(f11[1]) );
  CFD2QX1 \f03_reg[11]  ( .D(n283), .CP(clk), .CD(n887), .Q(f03[11]) );
  CFD2QX2 \f13_reg[21]  ( .D(n699), .CP(clk), .CD(n900), .Q(f13[21]) );
  CFD2QX1 \f17_reg[1]  ( .D(s17[1]), .CP(clk), .CD(n880), .Q(f17[1]) );
  CFD2QX1 \f21_reg[18]  ( .D(n619), .CP(clk), .CD(n911), .Q(f21[18]) );
  CFD2QX1 \f21_reg[21]  ( .D(n835), .CP(clk), .CD(n911), .Q(f21[21]) );
  CFD2QX2 \f12_reg[20]  ( .D(s12[20]), .CP(clk), .CD(n918), .Q(f12[20]) );
  CFD2QX2 \f02_reg[8]  ( .D(n774), .CP(clk), .CD(n897), .Q(f02[8]) );
  CFD2QX2 \f03_reg[8]  ( .D(n672), .CP(clk), .CD(n886), .Q(f03[8]) );
  CFD2QX1 \f23_reg[23]  ( .D(s23[23]), .CP(clk), .CD(n914), .Q(f23[23]) );
  CFD2QX1 \f14_reg[17]  ( .D(s14[17]), .CP(clk), .CD(n894), .Q(f14[17]) );
  CFD2QX2 \f13_reg[23]  ( .D(n714), .CP(clk), .CD(n900), .Q(f13[23]) );
  CFD2QX2 \f12_reg[24]  ( .D(s12[24]), .CP(clk), .CD(n919), .Q(f12[24]) );
  CFD2QX1 \f23_reg[14]  ( .D(s23[14]), .CP(clk), .CD(n913), .Q(f23[14]) );
  CNIVX1 U119 ( .A(n625), .Z(n119) );
  CNIVX3 U120 ( .A(f01[18]), .Z(n727) );
  CNIVXL U121 ( .A(f01[5]), .Z(n126) );
  CNIVXL U122 ( .A(f21[18]), .Z(n120) );
  CIVX1 U123 ( .A(f01[0]), .Z(n697) );
  CNIVX1 U124 ( .A(n698), .Z(n121) );
  CIVDX1 U125 ( .A(captC[11]), .Z1(n283) );
  CNIVX1 U126 ( .A(n825), .Z(n122) );
  CIVX2 U127 ( .A(n697), .Z(n698) );
  CDLY1XL U128 ( .A(f11[18]), .Z(n619) );
  CNIVX2 U129 ( .A(f12[19]), .Z(n828) );
  CNIVX1 U130 ( .A(f31[12]), .Z(n830) );
  CNIVX2 U131 ( .A(f01[1]), .Z(n684) );
  CNIVXL U132 ( .A(f01[15]), .Z(n833) );
  CNIVX1 U133 ( .A(f02[26]), .Z(n625) );
  CNIVXL U134 ( .A(f11[7]), .Z(n310) );
  CNIVX1 U135 ( .A(f02[14]), .Z(n705) );
  CNIVX1 U136 ( .A(f01[10]), .Z(n726) );
  CNIVX4 U137 ( .A(f12[2]), .Z(n123) );
  CNIVXL U138 ( .A(f02[15]), .Z(n124) );
  CNIVX1 U139 ( .A(f13[17]), .Z(n125) );
  CNIVX1 U140 ( .A(f01[13]), .Z(n127) );
  CNIVX1 U141 ( .A(f11[3]), .Z(n128) );
  CNIVX3 U142 ( .A(f11[6]), .Z(n130) );
  CNIVX1 U143 ( .A(n130), .Z(n129) );
  CNIVX3 U144 ( .A(f11[8]), .Z(n132) );
  CNIVX1 U145 ( .A(n132), .Z(n131) );
  CNIVX1 U146 ( .A(n134), .Z(n133) );
  CNIVX1 U147 ( .A(f11[10]), .Z(n134) );
  CDLY1XL U148 ( .A(f11[13]), .Z(n135) );
  CIVDX1 U149 ( .A(res_d[31]), .Z1(n137) );
  CNIVX1 U150 ( .A(n137), .Z(n136) );
  CIVDX1 U151 ( .A(res_d[30]), .Z1(n139) );
  CNIVX1 U152 ( .A(n139), .Z(n138) );
  CIVDX1 U153 ( .A(res_d[29]), .Z1(n141) );
  CNIVX1 U154 ( .A(n141), .Z(n140) );
  CIVDX1 U155 ( .A(res_d[28]), .Z1(n143) );
  CNIVX1 U156 ( .A(n143), .Z(n142) );
  CIVDX1 U157 ( .A(res_d[27]), .Z1(n145) );
  CNIVX1 U158 ( .A(n145), .Z(n144) );
  CIVDX1 U159 ( .A(res_d[26]), .Z1(n147) );
  CNIVX1 U160 ( .A(n147), .Z(n146) );
  CIVDX1 U161 ( .A(res_d[25]), .Z1(n149) );
  CNIVX1 U162 ( .A(n149), .Z(n148) );
  CIVDX1 U163 ( .A(res_d[24]), .Z1(n151) );
  CNIVX1 U164 ( .A(n151), .Z(n150) );
  CIVDX1 U165 ( .A(res_d[23]), .Z1(n153) );
  CNIVX1 U166 ( .A(n153), .Z(n152) );
  CIVDX1 U167 ( .A(res_d[22]), .Z1(n155) );
  CNIVX1 U168 ( .A(n155), .Z(n154) );
  CIVDX1 U169 ( .A(res_d[21]), .Z1(n157) );
  CNIVX1 U170 ( .A(n157), .Z(n156) );
  CIVDX1 U171 ( .A(res_d[20]), .Z1(n159) );
  CNIVX1 U172 ( .A(n159), .Z(n158) );
  CIVDX1 U173 ( .A(res_d[19]), .Z1(n161) );
  CNIVX1 U174 ( .A(n161), .Z(n160) );
  CIVDX1 U175 ( .A(res_d[18]), .Z1(n163) );
  CNIVX1 U176 ( .A(n163), .Z(n162) );
  CIVDX1 U177 ( .A(res_d[17]), .Z1(n165) );
  CNIVX1 U178 ( .A(n165), .Z(n164) );
  CIVDX1 U179 ( .A(res_d[16]), .Z1(n167) );
  CNIVX1 U180 ( .A(n167), .Z(n166) );
  CIVDX1 U181 ( .A(res_d[15]), .Z1(n169) );
  CNIVX1 U182 ( .A(n169), .Z(n168) );
  CIVDX1 U183 ( .A(res_d[14]), .Z1(n171) );
  CNIVX1 U184 ( .A(n171), .Z(n170) );
  CIVDX1 U185 ( .A(res_d[13]), .Z1(n173) );
  CNIVX1 U186 ( .A(n173), .Z(n172) );
  CIVDX1 U187 ( .A(res_d[12]), .Z1(n175) );
  CNIVX1 U188 ( .A(n175), .Z(n174) );
  CIVDX1 U189 ( .A(res_d[11]), .Z1(n177) );
  CNIVX1 U190 ( .A(n177), .Z(n176) );
  CIVDX1 U191 ( .A(res_d[10]), .Z1(n179) );
  CNIVX1 U192 ( .A(n179), .Z(n178) );
  CIVDX1 U193 ( .A(res_d[9]), .Z1(n181) );
  CNIVX1 U194 ( .A(n181), .Z(n180) );
  CIVDX1 U195 ( .A(res_d[8]), .Z1(n183) );
  CNIVX1 U196 ( .A(n183), .Z(n182) );
  CIVDX1 U197 ( .A(res_d[7]), .Z1(n185) );
  CNIVX1 U198 ( .A(n185), .Z(n184) );
  CIVDX1 U199 ( .A(res_d[6]), .Z1(n187) );
  CNIVX1 U200 ( .A(n187), .Z(n186) );
  CIVDX1 U201 ( .A(res_d[5]), .Z1(n189) );
  CNIVX1 U202 ( .A(n189), .Z(n188) );
  CIVDX1 U203 ( .A(res_d[4]), .Z1(n191) );
  CNIVX1 U204 ( .A(n191), .Z(n190) );
  CIVDX1 U205 ( .A(res_d[3]), .Z1(n193) );
  CNIVX1 U206 ( .A(n193), .Z(n192) );
  CIVDX1 U207 ( .A(res_d[2]), .Z1(n195) );
  CNIVX1 U208 ( .A(n195), .Z(n194) );
  CIVDX1 U209 ( .A(res_d[1]), .Z1(n197) );
  CNIVX1 U210 ( .A(n197), .Z(n196) );
  CIVDX1 U211 ( .A(res_d[0]), .Z1(n199) );
  CNIVX1 U212 ( .A(n199), .Z(n198) );
  CIVDX1 U213 ( .A(all_in7), .Z1(n201) );
  CNIVX1 U214 ( .A(n201), .Z(n200) );
  CIVDX1 U215 ( .A(f15[0]), .Z1(n203) );
  CNIVX1 U216 ( .A(n203), .Z(n202) );
  CIVDX1 U217 ( .A(f15[2]), .Z1(n205) );
  CNIVX1 U218 ( .A(n205), .Z(n204) );
  CIVDX1 U219 ( .A(f15[3]), .Z1(n207) );
  CNIVX1 U220 ( .A(n207), .Z(n206) );
  CIVDX1 U221 ( .A(f15[4]), .Z1(n209) );
  CNIVX1 U222 ( .A(n209), .Z(n208) );
  CIVDX1 U223 ( .A(f15[5]), .Z1(n211) );
  CNIVX1 U224 ( .A(n211), .Z(n210) );
  CIVDX1 U225 ( .A(f15[6]), .Z1(n213) );
  CNIVX1 U226 ( .A(n213), .Z(n212) );
  CIVDX1 U227 ( .A(f15[7]), .Z1(n215) );
  CNIVX1 U228 ( .A(n215), .Z(n214) );
  CIVDX1 U229 ( .A(f15[8]), .Z1(n217) );
  CNIVX1 U230 ( .A(n217), .Z(n216) );
  CIVDX1 U231 ( .A(f15[9]), .Z1(n219) );
  CNIVX1 U232 ( .A(n219), .Z(n218) );
  CIVDX1 U233 ( .A(f15[10]), .Z1(n221) );
  CNIVX1 U234 ( .A(n221), .Z(n220) );
  CIVDX1 U235 ( .A(f15[11]), .Z1(n223) );
  CNIVX1 U236 ( .A(n223), .Z(n222) );
  CIVDX1 U237 ( .A(f15[12]), .Z1(n225) );
  CNIVX1 U238 ( .A(n225), .Z(n224) );
  CIVDX1 U239 ( .A(f15[13]), .Z1(n227) );
  CNIVX1 U240 ( .A(n227), .Z(n226) );
  CIVDX1 U241 ( .A(f15[14]), .Z1(n229) );
  CNIVX1 U242 ( .A(n229), .Z(n228) );
  CIVDX1 U243 ( .A(f15[15]), .Z1(n231) );
  CNIVX1 U244 ( .A(n231), .Z(n230) );
  CIVDX1 U245 ( .A(f15[16]), .Z1(n233) );
  CNIVX1 U246 ( .A(n233), .Z(n232) );
  CIVDX1 U247 ( .A(f15[17]), .Z1(n235) );
  CNIVX1 U248 ( .A(n235), .Z(n234) );
  CIVDX1 U249 ( .A(f15[18]), .Z1(n237) );
  CNIVX1 U250 ( .A(n237), .Z(n236) );
  CIVDX1 U251 ( .A(f15[19]), .Z1(n239) );
  CNIVX1 U252 ( .A(n239), .Z(n238) );
  CIVDX1 U253 ( .A(f15[20]), .Z1(n241) );
  CNIVX1 U254 ( .A(n241), .Z(n240) );
  CIVDX1 U255 ( .A(f15[21]), .Z1(n243) );
  CNIVX1 U256 ( .A(n243), .Z(n242) );
  CIVDX1 U257 ( .A(f15[22]), .Z1(n245) );
  CNIVX1 U258 ( .A(n245), .Z(n244) );
  CIVDX1 U259 ( .A(f15[23]), .Z1(n247) );
  CNIVX1 U260 ( .A(n247), .Z(n246) );
  CIVDX1 U261 ( .A(f15[24]), .Z1(n249) );
  CNIVX1 U262 ( .A(n249), .Z(n248) );
  CIVDX1 U263 ( .A(f15[25]), .Z1(n251) );
  CNIVX1 U264 ( .A(n251), .Z(n250) );
  CIVDX1 U265 ( .A(f15[26]), .Z1(n253) );
  CNIVX1 U266 ( .A(n253), .Z(n252) );
  CIVDX1 U267 ( .A(f15[27]), .Z1(n255) );
  CNIVX1 U268 ( .A(n255), .Z(n254) );
  CIVDX1 U269 ( .A(f15[28]), .Z1(n257) );
  CNIVX1 U270 ( .A(n257), .Z(n256) );
  CIVDX1 U271 ( .A(f15[29]), .Z1(n259) );
  CNIVX1 U272 ( .A(n259), .Z(n258) );
  CIVDX1 U273 ( .A(f15[30]), .Z1(n261) );
  CNIVX1 U274 ( .A(n261), .Z(n260) );
  CIVDX1 U275 ( .A(f15[31]), .Z1(n263) );
  CNIVX1 U276 ( .A(n263), .Z(n262) );
  CNIVX3 U277 ( .A(f03[0]), .Z(n265) );
  CNIVX1 U278 ( .A(n265), .Z(n264) );
  CIVDX1 U279 ( .A(all_in6), .Z1(n267) );
  CNIVX1 U280 ( .A(n267), .Z(n266) );
  CIVDX1 U281 ( .A(all_in5), .Z1(n269) );
  CNIVX1 U282 ( .A(n269), .Z(n268) );
  CIVDX1 U283 ( .A(all_in4), .Z1(n271) );
  CNIVX1 U284 ( .A(n271), .Z(n270) );
  CIVDX1 U285 ( .A(all_in3), .Z1(n273) );
  CNIVX1 U286 ( .A(n273), .Z(n272) );
  CIVDX1 U287 ( .A(all_in2), .Z1(n275) );
  CNIVX1 U288 ( .A(n275), .Z(n274) );
  CIVDX1 U289 ( .A(all_in1), .Z1(n277) );
  CNIVX1 U290 ( .A(n277), .Z(n276) );
  CIVDX1 U291 ( .A(all_in), .Z1(n279) );
  CNIVX1 U292 ( .A(n279), .Z(n278) );
  CNIVX1 U293 ( .A(n281), .Z(n280) );
  CNIVX1 U294 ( .A(f21[21]), .Z(n281) );
  CIVDX1 U295 ( .A(captC[13]), .Z1(n282) );
  CNIVX1 U296 ( .A(f11[22]), .Z(n284) );
  CNIVXL U297 ( .A(captC[27]), .Z(n553) );
  CNIVX1 U298 ( .A(n553), .Z(n285) );
  CNIVX1 U299 ( .A(n287), .Z(n286) );
  CNIVX1 U300 ( .A(f11[23]), .Z(n287) );
  CNIVX1 U301 ( .A(f11[20]), .Z(n288) );
  CNIVX1 U302 ( .A(f21[23]), .Z(n289) );
  CNIVX1 U303 ( .A(n291), .Z(n290) );
  CNIVX1 U304 ( .A(f11[24]), .Z(n291) );
  CIVX4 U305 ( .A(n292), .Z(n293) );
  CIVXL U306 ( .A(f11[25]), .Z(n292) );
  CNIVX1 U307 ( .A(n295), .Z(n294) );
  CNIVX1 U308 ( .A(f11[26]), .Z(n295) );
  CNIVX1 U309 ( .A(f11[27]), .Z(n296) );
  CNIVXL U310 ( .A(captC[29]), .Z(n555) );
  CNIVX1 U311 ( .A(n555), .Z(n297) );
  CNIVX2 U312 ( .A(f01[28]), .Z(n298) );
  CNIVX1 U313 ( .A(f21[26]), .Z(n299) );
  CNIVX1 U314 ( .A(f21[27]), .Z(n300) );
  CNIVX1 U315 ( .A(f01[30]), .Z(n301) );
  CNIVXL U316 ( .A(captB[28]), .Z(n558) );
  CNIVX1 U317 ( .A(n558), .Z(n302) );
  CNIVXL U318 ( .A(captB[30]), .Z(n559) );
  CNIVX1 U319 ( .A(n559), .Z(n303) );
  CNIVXL U320 ( .A(captA[28]), .Z(n561) );
  CNIVX1 U321 ( .A(n561), .Z(n304) );
  CNIVXL U322 ( .A(captA[30]), .Z(n562) );
  CNIVX1 U323 ( .A(n562), .Z(n305) );
  CIVX3 U324 ( .A(n307), .Z(n308) );
  CNIVX1 U325 ( .A(n308), .Z(n306) );
  CIVXL U326 ( .A(f11[11]), .Z(n307) );
  CNIVX1 U327 ( .A(n310), .Z(n309) );
  CNIVX1 U328 ( .A(f02[30]), .Z(n311) );
  CNIVX1 U329 ( .A(f11[28]), .Z(n312) );
  CNIVX2 U330 ( .A(f21[28]), .Z(n313) );
  CNIVX2 U331 ( .A(f21[29]), .Z(n314) );
  CNIVXL U332 ( .A(captC[28]), .Z(n554) );
  CNIVX1 U333 ( .A(n554), .Z(n315) );
  CNIVX1 U334 ( .A(n317), .Z(n316) );
  CNIVX1 U335 ( .A(n318), .Z(n317) );
  CNIVX1 U336 ( .A(f11[5]), .Z(n318) );
  CNIVX1 U337 ( .A(n320), .Z(n319) );
  CNIVX1 U338 ( .A(n321), .Z(n320) );
  CNIVX1 U339 ( .A(f11[9]), .Z(n321) );
  CNIVXL U340 ( .A(f11[12]), .Z(n322) );
  CNIVXL U341 ( .A(f11[14]), .Z(n323) );
  CIVX4 U342 ( .A(n324), .Z(n325) );
  CIVXL U343 ( .A(f11[2]), .Z(n324) );
  CNIVX1 U344 ( .A(n327), .Z(n326) );
  CNIVX1 U345 ( .A(n328), .Z(n327) );
  CNIVX1 U346 ( .A(f11[4]), .Z(n328) );
  CNIVX1 U347 ( .A(f11[30]), .Z(n329) );
  CIVDX1 U348 ( .A(f43[2]), .Z1(n331) );
  CNIVX1 U349 ( .A(n331), .Z(n330) );
  CIVDX1 U350 ( .A(f43[6]), .Z1(n333) );
  CNIVX1 U351 ( .A(n333), .Z(n332) );
  CIVDX1 U352 ( .A(f32[2]), .Z1(n335) );
  CNIVX1 U353 ( .A(n335), .Z(n334) );
  CIVDX1 U354 ( .A(f32[5]), .Z1(n337) );
  CNIVX1 U355 ( .A(n337), .Z(n336) );
  CIVDX1 U356 ( .A(f32[6]), .Z1(n339) );
  CNIVX1 U357 ( .A(n339), .Z(n338) );
  CIVDX1 U358 ( .A(f25[2]), .Z1(n341) );
  CNIVX1 U359 ( .A(n341), .Z(n340) );
  CIVDX1 U360 ( .A(f25[6]), .Z1(n343) );
  CNIVX1 U361 ( .A(n343), .Z(n342) );
  CIVDX1 U362 ( .A(f43[12]), .Z1(n345) );
  CNIVX1 U363 ( .A(n345), .Z(n344) );
  CIVDX1 U364 ( .A(f43[13]), .Z1(n347) );
  CNIVX1 U365 ( .A(n347), .Z(n346) );
  CIVDX1 U366 ( .A(f43[14]), .Z1(n349) );
  CNIVX1 U367 ( .A(n349), .Z(n348) );
  CIVDX1 U368 ( .A(f43[15]), .Z1(n351) );
  CNIVX1 U369 ( .A(n351), .Z(n350) );
  CIVDX1 U370 ( .A(f32[12]), .Z1(n353) );
  CNIVX1 U371 ( .A(n353), .Z(n352) );
  CIVDX1 U372 ( .A(f32[13]), .Z1(n355) );
  CNIVX1 U373 ( .A(n355), .Z(n354) );
  CIVDX1 U374 ( .A(f32[14]), .Z1(n357) );
  CNIVX1 U375 ( .A(n357), .Z(n356) );
  CIVDX1 U376 ( .A(f32[15]), .Z1(n359) );
  CNIVX1 U377 ( .A(n359), .Z(n358) );
  CIVDX1 U378 ( .A(f43[0]), .Z1(n361) );
  CNIVX1 U379 ( .A(n361), .Z(n360) );
  CIVDX1 U380 ( .A(f43[4]), .Z1(n363) );
  CNIVX1 U381 ( .A(n363), .Z(n362) );
  CIVDX1 U382 ( .A(f43[5]), .Z1(n365) );
  CNIVX1 U383 ( .A(n365), .Z(n364) );
  CIVDX1 U384 ( .A(f43[7]), .Z1(n367) );
  CNIVX1 U385 ( .A(n367), .Z(n366) );
  CIVDX1 U386 ( .A(f43[8]), .Z1(n369) );
  CNIVX1 U387 ( .A(n369), .Z(n368) );
  CIVDX1 U388 ( .A(f43[9]), .Z1(n371) );
  CNIVX1 U389 ( .A(n371), .Z(n370) );
  CIVDX1 U390 ( .A(f43[10]), .Z1(n373) );
  CNIVX1 U391 ( .A(n373), .Z(n372) );
  CIVDX1 U392 ( .A(f43[11]), .Z1(n375) );
  CNIVX1 U393 ( .A(n375), .Z(n374) );
  CIVDX1 U394 ( .A(f32[0]), .Z1(n377) );
  CNIVX1 U395 ( .A(n377), .Z(n376) );
  CIVDX1 U396 ( .A(f32[4]), .Z1(n379) );
  CNIVX1 U397 ( .A(n379), .Z(n378) );
  CIVDX1 U398 ( .A(f32[7]), .Z1(n381) );
  CNIVX1 U399 ( .A(n381), .Z(n380) );
  CIVDX1 U400 ( .A(f32[8]), .Z1(n383) );
  CNIVX1 U401 ( .A(n383), .Z(n382) );
  CIVDX1 U402 ( .A(f32[9]), .Z1(n385) );
  CNIVX1 U403 ( .A(n385), .Z(n384) );
  CIVDX1 U404 ( .A(f32[10]), .Z1(n387) );
  CNIVX1 U405 ( .A(n387), .Z(n386) );
  CIVDX1 U406 ( .A(f32[11]), .Z1(n389) );
  CNIVX1 U407 ( .A(n389), .Z(n388) );
  CIVDX1 U408 ( .A(f25[0]), .Z1(n391) );
  CNIVX1 U409 ( .A(n391), .Z(n390) );
  CIVDX1 U410 ( .A(f25[4]), .Z1(n393) );
  CNIVX1 U411 ( .A(n393), .Z(n392) );
  CIVDX1 U412 ( .A(f25[5]), .Z1(n395) );
  CNIVX1 U413 ( .A(n395), .Z(n394) );
  CIVDX1 U414 ( .A(f25[7]), .Z1(n397) );
  CNIVX1 U415 ( .A(n397), .Z(n396) );
  CIVDX1 U416 ( .A(f25[8]), .Z1(n399) );
  CNIVX1 U417 ( .A(n399), .Z(n398) );
  CIVDX1 U418 ( .A(f25[9]), .Z1(n401) );
  CNIVX1 U419 ( .A(n401), .Z(n400) );
  CIVDX1 U420 ( .A(f25[10]), .Z1(n403) );
  CNIVX1 U421 ( .A(n403), .Z(n402) );
  CIVDX1 U422 ( .A(f25[11]), .Z1(n405) );
  CNIVX1 U423 ( .A(n405), .Z(n404) );
  CIVDX1 U424 ( .A(f25[12]), .Z1(n407) );
  CNIVX1 U425 ( .A(n407), .Z(n406) );
  CIVDX1 U426 ( .A(f25[13]), .Z1(n409) );
  CNIVX1 U427 ( .A(n409), .Z(n408) );
  CIVDX1 U428 ( .A(f25[14]), .Z1(n411) );
  CNIVX1 U429 ( .A(n411), .Z(n410) );
  CIVDX1 U430 ( .A(f25[15]), .Z1(n413) );
  CNIVX1 U431 ( .A(n413), .Z(n412) );
  CIVDX1 U432 ( .A(f43[1]), .Z1(n415) );
  CNIVX1 U433 ( .A(n415), .Z(n414) );
  CIVDX1 U434 ( .A(f43[3]), .Z1(n417) );
  CNIVX1 U435 ( .A(n417), .Z(n416) );
  CIVDX1 U436 ( .A(f32[1]), .Z1(n419) );
  CNIVX1 U437 ( .A(n419), .Z(n418) );
  CIVDX1 U438 ( .A(f32[3]), .Z1(n421) );
  CNIVX1 U439 ( .A(n421), .Z(n420) );
  CIVDX1 U440 ( .A(f25[3]), .Z1(n423) );
  CNIVX1 U441 ( .A(n423), .Z(n422) );
  CIVDX1 U442 ( .A(f43[16]), .Z1(n425) );
  CNIVX1 U443 ( .A(n425), .Z(n424) );
  CIVDX1 U444 ( .A(f43[17]), .Z1(n427) );
  CNIVX1 U445 ( .A(n427), .Z(n426) );
  CIVDX1 U446 ( .A(f43[18]), .Z1(n429) );
  CNIVX1 U447 ( .A(n429), .Z(n428) );
  CIVDX1 U448 ( .A(f32[16]), .Z1(n431) );
  CNIVX1 U449 ( .A(n431), .Z(n430) );
  CIVDX1 U450 ( .A(f32[17]), .Z1(n433) );
  CNIVX1 U451 ( .A(n433), .Z(n432) );
  CIVDX1 U452 ( .A(f32[18]), .Z1(n435) );
  CNIVX1 U453 ( .A(n435), .Z(n434) );
  CIVDX1 U454 ( .A(f32[19]), .Z1(n437) );
  CNIVX1 U455 ( .A(n437), .Z(n436) );
  CIVDX1 U456 ( .A(f25[16]), .Z1(n439) );
  CNIVX1 U457 ( .A(n439), .Z(n438) );
  CIVDX1 U458 ( .A(f25[17]), .Z1(n441) );
  CNIVX1 U459 ( .A(n441), .Z(n440) );
  CIVDX1 U460 ( .A(f25[18]), .Z1(n443) );
  CNIVX1 U461 ( .A(n443), .Z(n442) );
  CIVDX1 U462 ( .A(f25[19]), .Z1(n445) );
  CNIVX1 U463 ( .A(n445), .Z(n444) );
  CNIVXL U464 ( .A(captC[30]), .Z(n556) );
  CNIVX1 U465 ( .A(n556), .Z(n446) );
  CNIVX3 U466 ( .A(f01[4]), .Z(n447) );
  CNIVX1 U467 ( .A(n449), .Z(n448) );
  CNIVX1 U468 ( .A(f21[2]), .Z(n449) );
  CNIVX1 U469 ( .A(n451), .Z(n450) );
  CNIVX1 U470 ( .A(f21[3]), .Z(n451) );
  CNIVX1 U471 ( .A(n453), .Z(n452) );
  CNIVX1 U472 ( .A(f21[4]), .Z(n453) );
  CNIVX1 U473 ( .A(n455), .Z(n454) );
  CNIVX1 U474 ( .A(f21[5]), .Z(n455) );
  CNIVX1 U475 ( .A(n457), .Z(n456) );
  CNIVX1 U476 ( .A(f21[7]), .Z(n457) );
  CNIVX1 U477 ( .A(n459), .Z(n458) );
  CNIVX1 U478 ( .A(f21[6]), .Z(n459) );
  CNIVX1 U479 ( .A(n461), .Z(n460) );
  CNIVX1 U480 ( .A(f21[8]), .Z(n461) );
  CNIVX1 U481 ( .A(n463), .Z(n462) );
  CNIVX1 U482 ( .A(f21[9]), .Z(n463) );
  CIVX3 U483 ( .A(n464), .Z(n465) );
  CIVXL U484 ( .A(f21[11]), .Z(n464) );
  CNIVX1 U485 ( .A(n467), .Z(n466) );
  CNIVX1 U486 ( .A(f21[10]), .Z(n467) );
  CNIVX1 U487 ( .A(n469), .Z(n468) );
  CNIVX1 U488 ( .A(f21[12]), .Z(n469) );
  CNIVX1 U489 ( .A(n471), .Z(n470) );
  CNIVX1 U490 ( .A(f21[15]), .Z(n471) );
  CNIVX1 U491 ( .A(n473), .Z(n472) );
  CNIVX1 U492 ( .A(f21[30]), .Z(n473) );
  CNIVXL U493 ( .A(captB[31]), .Z(n560) );
  CNIVX1 U494 ( .A(n560), .Z(n474) );
  CNIVXL U495 ( .A(captA[31]), .Z(n563) );
  CNIVX1 U496 ( .A(n563), .Z(n475) );
  CIVDX1 U497 ( .A(f43[19]), .Z1(n477) );
  CNIVX1 U498 ( .A(n477), .Z(n476) );
  CIVDX1 U499 ( .A(f43[20]), .Z1(n479) );
  CNIVX1 U500 ( .A(n479), .Z(n478) );
  CIVDX1 U501 ( .A(f43[21]), .Z1(n481) );
  CNIVX1 U502 ( .A(n481), .Z(n480) );
  CIVDX1 U503 ( .A(f43[22]), .Z1(n483) );
  CNIVX1 U504 ( .A(n483), .Z(n482) );
  CIVDX1 U505 ( .A(f43[23]), .Z1(n485) );
  CNIVX1 U506 ( .A(n485), .Z(n484) );
  CIVDX1 U507 ( .A(f43[24]), .Z1(n487) );
  CNIVX1 U508 ( .A(n487), .Z(n486) );
  CIVDX1 U509 ( .A(f43[25]), .Z1(n489) );
  CNIVX1 U510 ( .A(n489), .Z(n488) );
  CIVDX1 U511 ( .A(f43[26]), .Z1(n491) );
  CNIVX1 U512 ( .A(n491), .Z(n490) );
  CIVDX1 U513 ( .A(f43[27]), .Z1(n493) );
  CNIVX1 U514 ( .A(n493), .Z(n492) );
  CIVDX1 U515 ( .A(f32[20]), .Z1(n495) );
  CNIVX1 U516 ( .A(n495), .Z(n494) );
  CIVDX1 U517 ( .A(f32[21]), .Z1(n497) );
  CNIVX1 U518 ( .A(n497), .Z(n496) );
  CIVDX1 U519 ( .A(f32[22]), .Z1(n499) );
  CNIVX1 U520 ( .A(n499), .Z(n498) );
  CIVDX1 U521 ( .A(f32[23]), .Z1(n501) );
  CNIVX1 U522 ( .A(n501), .Z(n500) );
  CIVDX1 U523 ( .A(f32[24]), .Z1(n503) );
  CNIVX1 U524 ( .A(n503), .Z(n502) );
  CIVDX1 U525 ( .A(f32[25]), .Z1(n505) );
  CNIVX1 U526 ( .A(n505), .Z(n504) );
  CIVDX1 U527 ( .A(f32[26]), .Z1(n507) );
  CNIVX1 U528 ( .A(n507), .Z(n506) );
  CIVDX1 U529 ( .A(f32[27]), .Z1(n509) );
  CNIVX1 U530 ( .A(n509), .Z(n508) );
  CIVDX1 U531 ( .A(f25[20]), .Z1(n511) );
  CNIVX1 U532 ( .A(n511), .Z(n510) );
  CIVDX1 U533 ( .A(f25[21]), .Z1(n513) );
  CNIVX1 U534 ( .A(n513), .Z(n512) );
  CIVDX1 U535 ( .A(f25[22]), .Z1(n515) );
  CNIVX1 U536 ( .A(n515), .Z(n514) );
  CIVDX1 U537 ( .A(f25[23]), .Z1(n517) );
  CNIVX1 U538 ( .A(n517), .Z(n516) );
  CIVDX1 U539 ( .A(f25[24]), .Z1(n519) );
  CNIVX1 U540 ( .A(n519), .Z(n518) );
  CIVDX1 U541 ( .A(f25[25]), .Z1(n521) );
  CNIVX1 U542 ( .A(n521), .Z(n520) );
  CIVDX1 U543 ( .A(f25[26]), .Z1(n523) );
  CNIVX1 U544 ( .A(n523), .Z(n522) );
  CIVDX1 U545 ( .A(f25[27]), .Z1(n525) );
  CNIVX1 U546 ( .A(n525), .Z(n524) );
  CNIVXL U547 ( .A(captC[31]), .Z(n557) );
  CNIVX1 U548 ( .A(n557), .Z(n526) );
  CNIVX1 U549 ( .A(n528), .Z(n527) );
  CNIVX1 U550 ( .A(f21[31]), .Z(n528) );
  CIVDX1 U551 ( .A(f43[31]), .Z1(n530) );
  CNIVX1 U552 ( .A(n530), .Z(n529) );
  CIVDX1 U553 ( .A(f32[31]), .Z1(n532) );
  CNIVX1 U554 ( .A(n532), .Z(n531) );
  CIVDX1 U555 ( .A(f25[31]), .Z1(n534) );
  CNIVX1 U556 ( .A(n534), .Z(n533) );
  CIVDX1 U557 ( .A(f43[28]), .Z1(n536) );
  CNIVX1 U558 ( .A(n536), .Z(n535) );
  CIVDX1 U559 ( .A(f43[29]), .Z1(n538) );
  CNIVX1 U560 ( .A(n538), .Z(n537) );
  CIVDX1 U561 ( .A(f43[30]), .Z1(n540) );
  CNIVX1 U562 ( .A(n540), .Z(n539) );
  CIVDX1 U563 ( .A(f32[28]), .Z1(n542) );
  CNIVX1 U564 ( .A(n542), .Z(n541) );
  CIVDX1 U565 ( .A(f32[29]), .Z1(n544) );
  CNIVX1 U566 ( .A(n544), .Z(n543) );
  CIVDX1 U567 ( .A(f32[30]), .Z1(n546) );
  CNIVX1 U568 ( .A(n546), .Z(n545) );
  CIVDX1 U569 ( .A(f25[28]), .Z1(n548) );
  CNIVX1 U570 ( .A(n548), .Z(n547) );
  CIVDX1 U571 ( .A(f25[29]), .Z1(n550) );
  CNIVX1 U572 ( .A(n550), .Z(n549) );
  CIVDX1 U573 ( .A(f25[30]), .Z1(n552) );
  CNIVX1 U574 ( .A(n552), .Z(n551) );
  CNIVX1 U575 ( .A(n565), .Z(n564) );
  CNIVX1 U576 ( .A(f11[0]), .Z(n565) );
  CNIVX1 U577 ( .A(n567), .Z(n566) );
  CNIVX1 U578 ( .A(f11[17]), .Z(n567) );
  CNIVX1 U579 ( .A(n569), .Z(n568) );
  CNIVX1 U580 ( .A(n570), .Z(n569) );
  CNIVX1 U581 ( .A(f02[17]), .Z(n570) );
  CIVDX1 U582 ( .A(captB[21]), .Z1(n571) );
  CNIVX3 U583 ( .A(f02[29]), .Z(n572) );
  CIVDX1 U584 ( .A(captA[19]), .Z1(n573) );
  CIVDX1 U585 ( .A(captA[5]), .Z1(n574) );
  CNIVX1 U586 ( .A(n576), .Z(n575) );
  CNIVX1 U587 ( .A(f02[1]), .Z(n576) );
  CNIVX1 U588 ( .A(n578), .Z(n577) );
  CNIVX1 U589 ( .A(captC[4]), .Z(n578) );
  CIVDX1 U590 ( .A(captA[13]), .Z1(n579) );
  CNIVX1 U591 ( .A(n581), .Z(n580) );
  CNIVX1 U592 ( .A(captC[5]), .Z(n581) );
  CNIVX1 U593 ( .A(n583), .Z(n582) );
  CNIVX1 U594 ( .A(f02[7]), .Z(n583) );
  CNIVX1 U595 ( .A(n585), .Z(n584) );
  CNIVX1 U596 ( .A(f02[3]), .Z(n585) );
  CNIVX1 U597 ( .A(n587), .Z(n586) );
  CNIVX1 U598 ( .A(f02[11]), .Z(n587) );
  CNIVXL U599 ( .A(f01[12]), .Z(n588) );
  CNIVX1 U600 ( .A(n590), .Z(n589) );
  CNIVX1 U601 ( .A(f01[11]), .Z(n590) );
  CNIVX1 U602 ( .A(n592), .Z(n591) );
  CNIVX1 U603 ( .A(f02[13]), .Z(n592) );
  CNIVX1 U604 ( .A(n127), .Z(n593) );
  CNIVX1 U605 ( .A(n595), .Z(n594) );
  CNIVX1 U606 ( .A(captC[15]), .Z(n595) );
  CNIVX1 U607 ( .A(n597), .Z(n596) );
  CNIVX1 U608 ( .A(n128), .Z(n597) );
  CNIVX1 U609 ( .A(n599), .Z(n598) );
  CNIVX1 U610 ( .A(captC[9]), .Z(n599) );
  CNIVX1 U611 ( .A(n601), .Z(n600) );
  CNIVX1 U612 ( .A(f02[5]), .Z(n601) );
  CNIVX1 U613 ( .A(n603), .Z(n602) );
  CNIVX1 U614 ( .A(captB[25]), .Z(n603) );
  CNIVX1 U615 ( .A(n605), .Z(n604) );
  CNIVX1 U616 ( .A(f01[26]), .Z(n605) );
  CNIVX3 U617 ( .A(f01[16]), .Z(n606) );
  CIVDX1 U618 ( .A(captB[19]), .Z1(n607) );
  CNIVX1 U619 ( .A(n609), .Z(n608) );
  CNIVX1 U620 ( .A(n610), .Z(n609) );
  CNIVX1 U621 ( .A(f02[19]), .Z(n610) );
  CIVDX1 U622 ( .A(captA[16]), .Z1(n611) );
  CNIVX1 U623 ( .A(n613), .Z(n612) );
  CNIVX1 U624 ( .A(f02[9]), .Z(n613) );
  CNIVX1 U625 ( .A(f11[16]), .Z(n614) );
  CNIVX1 U626 ( .A(n616), .Z(n615) );
  CNIVX1 U627 ( .A(captC[16]), .Z(n616) );
  CIVDX1 U628 ( .A(captA[26]), .Z1(n617) );
  CNIVX1 U629 ( .A(f21[16]), .Z(n618) );
  CNIVX1 U630 ( .A(n621), .Z(n620) );
  CNIVX1 U631 ( .A(captB[23]), .Z(n621) );
  CNIVX1 U632 ( .A(n623), .Z(n622) );
  CNIVX1 U633 ( .A(f01[6]), .Z(n623) );
  CIVDX1 U634 ( .A(captA[15]), .Z1(n624) );
  CIVDX1 U635 ( .A(captB[26]), .Z1(n626) );
  CNIVX3 U636 ( .A(f02[10]), .Z(n627) );
  CIVDX1 U637 ( .A(captB[6]), .Z1(n628) );
  CIVDX1 U638 ( .A(captA[22]), .Z1(n629) );
  CNIVX1 U639 ( .A(n631), .Z(n630) );
  CNIVX1 U640 ( .A(f01[14]), .Z(n631) );
  CNIVX1 U641 ( .A(n633), .Z(n632) );
  CNIVX1 U642 ( .A(captA[12]), .Z(n633) );
  CNIVXL U643 ( .A(f02[6]), .Z(n634) );
  CIVDX1 U644 ( .A(captB[17]), .Z1(n635) );
  CIVDX1 U645 ( .A(captB[9]), .Z1(n636) );
  CIVDX1 U646 ( .A(captA[20]), .Z1(n637) );
  CIVDX1 U647 ( .A(captA[29]), .Z1(n638) );
  CIVDX1 U648 ( .A(captB[29]), .Z1(n639) );
  CNIVX1 U649 ( .A(f02[28]), .Z(n640) );
  CIVDX1 U650 ( .A(captC[23]), .Z1(n641) );
  CNIVX1 U651 ( .A(n643), .Z(n642) );
  CNIVX1 U652 ( .A(n644), .Z(n643) );
  CNIVX1 U653 ( .A(f01[23]), .Z(n644) );
  CIVXL U654 ( .A(n834), .Z(n835) );
  CNIVX1 U655 ( .A(n646), .Z(n645) );
  CNIVX1 U656 ( .A(captA[6]), .Z(n646) );
  CIVDX1 U657 ( .A(captA[14]), .Z1(n647) );
  CNIVX1 U658 ( .A(n649), .Z(n648) );
  CNIVX1 U659 ( .A(captB[10]), .Z(n649) );
  CNIVX1 U660 ( .A(n126), .Z(n650) );
  CNIVX1 U661 ( .A(n652), .Z(n651) );
  CNIVX1 U662 ( .A(n653), .Z(n652) );
  CNIVX1 U663 ( .A(f01[21]), .Z(n653) );
  CIVDX1 U664 ( .A(captA[21]), .Z1(n654) );
  CNIVX3 U665 ( .A(f01[25]), .Z(n656) );
  CNIVX1 U666 ( .A(n656), .Z(n655) );
  CNIVX1 U667 ( .A(n658), .Z(n657) );
  CNIVX1 U668 ( .A(captA[25]), .Z(n658) );
  CNIVX1 U669 ( .A(n660), .Z(n659) );
  CNIVX1 U670 ( .A(f21[1]), .Z(n660) );
  CDLY1XL U671 ( .A(f21[13]), .Z(n661) );
  CNIVX1 U672 ( .A(n663), .Z(n662) );
  CNIVX1 U673 ( .A(f21[14]), .Z(n663) );
  CNIVX3 U674 ( .A(f01[29]), .Z(n664) );
  CNIVX1 U675 ( .A(n666), .Z(n665) );
  CNIVX1 U676 ( .A(f01[19]), .Z(n666) );
  CIVDX1 U677 ( .A(captC[26]), .Z1(n667) );
  CNIVX1 U678 ( .A(n669), .Z(n668) );
  CNIVX1 U679 ( .A(f01[7]), .Z(n669) );
  CNIVXL U680 ( .A(captC[25]), .Z(n671) );
  CNIVX1 U681 ( .A(n671), .Z(n670) );
  CNIVX1 U682 ( .A(n673), .Z(n672) );
  CNIVX1 U683 ( .A(captC[8]), .Z(n673) );
  CIVDX1 U684 ( .A(captB[22]), .Z1(n674) );
  CNIVX1 U685 ( .A(n676), .Z(n675) );
  CNIVX1 U686 ( .A(n677), .Z(n676) );
  CNIVX1 U687 ( .A(f01[22]), .Z(n677) );
  CNIVX1 U688 ( .A(n679), .Z(n678) );
  CNIVX1 U689 ( .A(n680), .Z(n679) );
  CNIVX1 U690 ( .A(f01[17]), .Z(n680) );
  CIVDX1 U691 ( .A(captA[24]), .Z1(n681) );
  CIVDX1 U692 ( .A(captA[17]), .Z1(n682) );
  CNIVX1 U693 ( .A(n684), .Z(n683) );
  CNIVX1 U694 ( .A(n686), .Z(n685) );
  CNIVX1 U695 ( .A(captA[23]), .Z(n686) );
  CNIVX1 U696 ( .A(f21[17]), .Z(n687) );
  CNIVX1 U697 ( .A(n689), .Z(n688) );
  CNIVX1 U698 ( .A(n690), .Z(n689) );
  CNIVX1 U699 ( .A(f11[1]), .Z(n690) );
  CNIVX1 U700 ( .A(n692), .Z(n691) );
  CNIVX1 U701 ( .A(f01[3]), .Z(n692) );
  CNIVXL U702 ( .A(f02[0]), .Z(n693) );
  CNIVX1 U703 ( .A(n695), .Z(n694) );
  CNIVX1 U704 ( .A(f02[4]), .Z(n695) );
  CNIVX1 U705 ( .A(n698), .Z(n696) );
  CNIVX1 U706 ( .A(n700), .Z(n699) );
  CNIVX1 U707 ( .A(n701), .Z(n700) );
  CNIVX1 U708 ( .A(f02[21]), .Z(n701) );
  CNIVXL U709 ( .A(f02[2]), .Z(n702) );
  CNIVX1 U710 ( .A(n704), .Z(n703) );
  CNIVX1 U711 ( .A(f02[12]), .Z(n704) );
  CNIVX1 U712 ( .A(n707), .Z(n706) );
  CNIVX1 U713 ( .A(f02[16]), .Z(n707) );
  CNIVX1 U714 ( .A(n709), .Z(n708) );
  CNIVX1 U715 ( .A(f02[18]), .Z(n709) );
  CNIVX1 U716 ( .A(n711), .Z(n710) );
  CNIVX1 U717 ( .A(f02[20]), .Z(n711) );
  CNIVX1 U718 ( .A(n713), .Z(n712) );
  CNIVX1 U719 ( .A(f02[22]), .Z(n713) );
  CNIVX1 U720 ( .A(n715), .Z(n714) );
  CNIVX1 U721 ( .A(n716), .Z(n715) );
  CNIVX1 U722 ( .A(f02[23]), .Z(n716) );
  CNIVX1 U723 ( .A(n718), .Z(n717) );
  CNIVX1 U724 ( .A(f02[24]), .Z(n718) );
  CNIVX1 U725 ( .A(n720), .Z(n719) );
  CNIVX1 U726 ( .A(n721), .Z(n720) );
  CNIVX1 U727 ( .A(f02[25]), .Z(n721) );
  CNIVX1 U728 ( .A(f02[27]), .Z(n722) );
  CIVDX1 U729 ( .A(captC[24]), .Z1(n723) );
  CNIVX1 U730 ( .A(n725), .Z(n724) );
  CNIVX1 U731 ( .A(f01[2]), .Z(n725) );
  CNIVX3 U732 ( .A(f01[20]), .Z(n728) );
  CNIVX1 U733 ( .A(n730), .Z(n729) );
  CNIVX1 U734 ( .A(f01[24]), .Z(n730) );
  CNIVX1 U735 ( .A(f01[27]), .Z(n731) );
  CNIVX1 U736 ( .A(n733), .Z(n732) );
  CNIVX1 U737 ( .A(captC[0]), .Z(n733) );
  CNIVX1 U738 ( .A(n735), .Z(n734) );
  CNIVX1 U739 ( .A(captC[1]), .Z(n735) );
  CNIVX1 U740 ( .A(n737), .Z(n736) );
  CNIVX1 U741 ( .A(captC[2]), .Z(n737) );
  CNIVX1 U742 ( .A(n739), .Z(n738) );
  CNIVX1 U743 ( .A(captC[3]), .Z(n739) );
  CNIVX1 U744 ( .A(n741), .Z(n740) );
  CNIVX1 U745 ( .A(captC[6]), .Z(n741) );
  CNIVX1 U746 ( .A(n743), .Z(n742) );
  CNIVX1 U747 ( .A(captC[10]), .Z(n743) );
  CNIVX1 U748 ( .A(n745), .Z(n744) );
  CNIVX1 U749 ( .A(captC[12]), .Z(n745) );
  CNIVX1 U750 ( .A(n747), .Z(n746) );
  CNIVX1 U751 ( .A(captC[14]), .Z(n747) );
  CNIVX1 U752 ( .A(n749), .Z(n748) );
  CNIVX1 U753 ( .A(captC[17]), .Z(n749) );
  CNIVX1 U754 ( .A(n751), .Z(n750) );
  CNIVX1 U755 ( .A(captC[18]), .Z(n751) );
  CNIVX1 U756 ( .A(n753), .Z(n752) );
  CNIVX1 U757 ( .A(captC[19]), .Z(n753) );
  CNIVX1 U758 ( .A(n755), .Z(n754) );
  CNIVX1 U759 ( .A(captC[20]), .Z(n755) );
  CNIVX1 U760 ( .A(n757), .Z(n756) );
  CNIVX1 U761 ( .A(captC[21]), .Z(n757) );
  CNIVX1 U762 ( .A(n759), .Z(n758) );
  CNIVX1 U763 ( .A(captC[22]), .Z(n759) );
  CNIVX1 U764 ( .A(n761), .Z(n760) );
  CNIVX1 U765 ( .A(captB[0]), .Z(n761) );
  CNIVX1 U766 ( .A(n763), .Z(n762) );
  CNIVX1 U767 ( .A(captB[1]), .Z(n763) );
  CNIVX1 U768 ( .A(n765), .Z(n764) );
  CNIVX1 U769 ( .A(captB[2]), .Z(n765) );
  CNIVX1 U770 ( .A(n767), .Z(n766) );
  CNIVX1 U771 ( .A(captB[3]), .Z(n767) );
  CNIVX1 U772 ( .A(n769), .Z(n768) );
  CNIVX1 U773 ( .A(captB[4]), .Z(n769) );
  CNIVX1 U774 ( .A(n771), .Z(n770) );
  CNIVX1 U775 ( .A(captB[5]), .Z(n771) );
  CNIVX1 U776 ( .A(n773), .Z(n772) );
  CNIVX1 U777 ( .A(captB[7]), .Z(n773) );
  CNIVX1 U778 ( .A(n775), .Z(n774) );
  CNIVX1 U779 ( .A(captB[8]), .Z(n775) );
  CNIVX1 U780 ( .A(n777), .Z(n776) );
  CNIVX1 U781 ( .A(captB[11]), .Z(n777) );
  CNIVX1 U782 ( .A(n779), .Z(n778) );
  CNIVX1 U783 ( .A(captB[12]), .Z(n779) );
  CNIVX1 U784 ( .A(n781), .Z(n780) );
  CNIVX1 U785 ( .A(captB[13]), .Z(n781) );
  CNIVX1 U786 ( .A(n783), .Z(n782) );
  CNIVX1 U787 ( .A(captB[14]), .Z(n783) );
  CNIVX1 U788 ( .A(n785), .Z(n784) );
  CNIVX1 U789 ( .A(captB[15]), .Z(n785) );
  CNIVX1 U790 ( .A(n787), .Z(n786) );
  CNIVX1 U791 ( .A(captB[16]), .Z(n787) );
  CNIVX1 U792 ( .A(n789), .Z(n788) );
  CNIVX1 U793 ( .A(captB[18]), .Z(n789) );
  CNIVX1 U794 ( .A(n791), .Z(n790) );
  CNIVX1 U795 ( .A(f01[9]), .Z(n791) );
  CNIVX1 U796 ( .A(n793), .Z(n792) );
  CNIVX1 U797 ( .A(captB[27]), .Z(n793) );
  CNIVX1 U798 ( .A(n795), .Z(n794) );
  CNIVX1 U799 ( .A(captA[0]), .Z(n795) );
  CNIVX1 U800 ( .A(n797), .Z(n796) );
  CNIVX1 U801 ( .A(captA[1]), .Z(n797) );
  CNIVX1 U802 ( .A(n799), .Z(n798) );
  CNIVX1 U803 ( .A(captA[2]), .Z(n799) );
  CNIVX1 U804 ( .A(n801), .Z(n800) );
  CNIVX1 U805 ( .A(captA[3]), .Z(n801) );
  CNIVX1 U806 ( .A(n803), .Z(n802) );
  CNIVX1 U807 ( .A(captA[4]), .Z(n803) );
  CNIVX1 U808 ( .A(n805), .Z(n804) );
  CNIVX1 U809 ( .A(captA[7]), .Z(n805) );
  CNIVX1 U810 ( .A(n807), .Z(n806) );
  CNIVX1 U811 ( .A(captA[8]), .Z(n807) );
  CNIVX1 U812 ( .A(n809), .Z(n808) );
  CNIVX1 U813 ( .A(captA[9]), .Z(n809) );
  CNIVX1 U814 ( .A(n811), .Z(n810) );
  CNIVX1 U815 ( .A(captA[10]), .Z(n811) );
  CNIVX1 U816 ( .A(n813), .Z(n812) );
  CNIVX1 U817 ( .A(captA[11]), .Z(n813) );
  CNIVX1 U818 ( .A(n815), .Z(n814) );
  CNIVX1 U819 ( .A(n816), .Z(n815) );
  CNIVX1 U820 ( .A(f21[0]), .Z(n816) );
  CNIVX1 U821 ( .A(n818), .Z(n817) );
  CNIVX1 U822 ( .A(captC[7]), .Z(n818) );
  CNIVX1 U823 ( .A(n820), .Z(n819) );
  CNIVX1 U824 ( .A(captA[27]), .Z(n820) );
  CNIVX3 U825 ( .A(f21[19]), .Z(n821) );
  CIVDX1 U826 ( .A(captA[18]), .Z1(n822) );
  CIVDX1 U827 ( .A(captB[24]), .Z1(n823) );
  CIVDX1 U828 ( .A(captB[20]), .Z1(n824) );
  CNIVXL U829 ( .A(f02[8]), .Z(n825) );
  CNIVX1 U830 ( .A(n827), .Z(n826) );
  CNIVX1 U831 ( .A(f01[8]), .Z(n827) );
  CNIVX1 U832 ( .A(f11[19]), .Z(n829) );
  CNR3XL U833 ( .A(n15), .B(n13), .C(n14), .Z(N6) );
  CNR2X1 U834 ( .A(N6), .B(n14), .Z(seen_d[1]) );
  CNR2X1 U835 ( .A(N6), .B(n13), .Z(seen_d[2]) );
  CNR2X1 U836 ( .A(N6), .B(n15), .Z(seen_d[0]) );
  CNIVX1 U837 ( .A(n926), .Z(n886) );
  CNIVX1 U838 ( .A(n926), .Z(n887) );
  CNIVX1 U839 ( .A(n926), .Z(n916) );
  CNIVX1 U840 ( .A(n926), .Z(n919) );
  CNIVX1 U841 ( .A(n926), .Z(n915) );
  CNIVX1 U842 ( .A(n926), .Z(n896) );
  CNIVX1 U843 ( .A(n926), .Z(n846) );
  CNIVX1 U844 ( .A(n926), .Z(n847) );
  CNIVX1 U845 ( .A(n926), .Z(n848) );
  CNIVX1 U846 ( .A(n926), .Z(n849) );
  CNIVX1 U847 ( .A(n926), .Z(n850) );
  CNIVX1 U848 ( .A(n926), .Z(n851) );
  CNIVX1 U849 ( .A(n926), .Z(n852) );
  CNIVX1 U850 ( .A(n926), .Z(n853) );
  CNIVX1 U851 ( .A(n926), .Z(n854) );
  CNIVX1 U852 ( .A(n926), .Z(n872) );
  CNIVX1 U853 ( .A(n926), .Z(n871) );
  CNIVX1 U854 ( .A(n926), .Z(n903) );
  CNIVX1 U855 ( .A(n926), .Z(n904) );
  CNIVX1 U856 ( .A(n926), .Z(n864) );
  CNIVX1 U857 ( .A(n926), .Z(n873) );
  CNIVX1 U858 ( .A(n926), .Z(n874) );
  CNIVX1 U859 ( .A(n926), .Z(n875) );
  CNIVX1 U860 ( .A(n926), .Z(n876) );
  CNIVX1 U861 ( .A(n926), .Z(n877) );
  CNIVX1 U862 ( .A(n926), .Z(n905) );
  CNIVX1 U863 ( .A(n926), .Z(n878) );
  CNIVX1 U864 ( .A(n926), .Z(n879) );
  CNIVX1 U865 ( .A(n926), .Z(n891) );
  CNIVX1 U866 ( .A(n926), .Z(n855) );
  CNIVX1 U867 ( .A(n926), .Z(n869) );
  CNIVX1 U868 ( .A(n926), .Z(n870) );
  CNIVX1 U869 ( .A(n926), .Z(n865) );
  CNIVX1 U870 ( .A(n926), .Z(n866) );
  CNIVX1 U871 ( .A(n926), .Z(n867) );
  CNIVX1 U872 ( .A(n926), .Z(n868) );
  CNIVX1 U873 ( .A(n926), .Z(n880) );
  CNIVX1 U874 ( .A(n926), .Z(n881) );
  CNIVX1 U875 ( .A(n926), .Z(n882) );
  CNIVX1 U876 ( .A(n926), .Z(n883) );
  CNIVX1 U877 ( .A(n926), .Z(n884) );
  CNIVX1 U878 ( .A(n926), .Z(n857) );
  CNIVX1 U879 ( .A(n926), .Z(n858) );
  CNIVX1 U880 ( .A(n926), .Z(n859) );
  CNIVX1 U881 ( .A(n926), .Z(n860) );
  CNIVX1 U882 ( .A(n926), .Z(n861) );
  CNIVX1 U883 ( .A(n926), .Z(n863) );
  CNIVX1 U884 ( .A(n926), .Z(n893) );
  CNIVX1 U885 ( .A(n926), .Z(n894) );
  CNIVX1 U886 ( .A(n926), .Z(n914) );
  CNIVX1 U887 ( .A(n926), .Z(n885) );
  CNIVX1 U888 ( .A(n926), .Z(n888) );
  CNIVX1 U889 ( .A(n926), .Z(n889) );
  CNIVX1 U890 ( .A(n926), .Z(n890) );
  CNIVX1 U891 ( .A(n926), .Z(n901) );
  CNIVX1 U892 ( .A(n926), .Z(n902) );
  CNIVX1 U893 ( .A(n926), .Z(n920) );
  CNIVX1 U894 ( .A(n926), .Z(n923) );
  CNIVX1 U895 ( .A(n926), .Z(n924) );
  CNIVX1 U896 ( .A(n926), .Z(n906) );
  CNIVX1 U897 ( .A(n926), .Z(n907) );
  CNIVX1 U898 ( .A(n926), .Z(n912) );
  CNIVX1 U899 ( .A(n926), .Z(n918) );
  CNIVX1 U900 ( .A(n926), .Z(n899) );
  CNIVX1 U901 ( .A(n926), .Z(n900) );
  CNIVX1 U902 ( .A(n926), .Z(n921) );
  CNIVX1 U903 ( .A(n926), .Z(n922) );
  CNIVX1 U904 ( .A(n926), .Z(n908) );
  CNIVX1 U905 ( .A(n926), .Z(n895) );
  CNIVX1 U906 ( .A(n926), .Z(n897) );
  CNIVX1 U907 ( .A(n926), .Z(n898) );
  CNIVX1 U908 ( .A(n926), .Z(n913) );
  CNIVX1 U909 ( .A(n926), .Z(n909) );
  CNIVX1 U910 ( .A(n926), .Z(n862) );
  CNIVX1 U911 ( .A(n926), .Z(n910) );
  CNIVX1 U912 ( .A(n926), .Z(n911) );
  CNIVX1 U913 ( .A(n926), .Z(n892) );
  CNIVX1 U914 ( .A(n926), .Z(n917) );
  CNIVX1 U915 ( .A(n926), .Z(n856) );
  CNIVX1 U916 ( .A(n926), .Z(n925) );
  CNR2IX1 U917 ( .B(pushC), .A(stopC), .Z(n845) );
  CNR2IX1 U918 ( .B(pushC), .A(stopC), .Z(n844) );
  CNR2IX1 U919 ( .B(pushB), .A(stopB), .Z(n843) );
  CNR2IX1 U920 ( .B(pushB), .A(stopB), .Z(n842) );
  CNR2IX1 U921 ( .B(pushA), .A(stopA), .Z(n841) );
  CNR2IX1 U922 ( .B(pushA), .A(stopA), .Z(n840) );
  CNR2IX1 U923 ( .B(pushC), .A(stopC), .Z(n16) );
  CNR2IX1 U924 ( .B(pushB), .A(stopB), .Z(n18) );
  CNR2IX1 U925 ( .B(pushA), .A(stopA), .Z(n20) );
  CNR2X1 U926 ( .A(stopB), .B(pushB), .Z(n14) );
  CNR2X1 U927 ( .A(pushA), .B(stopA), .Z(n13) );
  CNR2X1 U928 ( .A(pushC), .B(stopC), .Z(n15) );
  CIVX2 U929 ( .A(rst), .Z(n926) );
  CIVXL U933 ( .A(f13[19]), .Z(n831) );
  CIVX2 U934 ( .A(n831), .Z(n832) );
  CIVXL U935 ( .A(f11[21]), .Z(n834) );
  CIVXL U936 ( .A(f13[5]), .Z(n836) );
  CIVXL U937 ( .A(n836), .Z(n837) );
  CIVXL U938 ( .A(f13[3]), .Z(n838) );
  CIVXL U939 ( .A(n838), .Z(n839) );
  CMX2X1 U940 ( .A0(n563), .A1(A[31]), .S(n840), .Z(n117) );
  CMX2X1 U941 ( .A0(n562), .A1(A[30]), .S(n841), .Z(n116) );
  CMX2X1 U942 ( .A0(captA[29]), .A1(A[29]), .S(n20), .Z(n115) );
  CMX2X1 U943 ( .A0(n561), .A1(A[28]), .S(n840), .Z(n114) );
  CMX2X1 U944 ( .A0(captA[27]), .A1(A[27]), .S(n841), .Z(n113) );
  CMX2X1 U945 ( .A0(captA[26]), .A1(A[26]), .S(n20), .Z(n112) );
  CMX2X1 U946 ( .A0(captA[25]), .A1(A[25]), .S(n840), .Z(n111) );
  CMX2X1 U947 ( .A0(captA[24]), .A1(A[24]), .S(n841), .Z(n110) );
  CMX2X1 U948 ( .A0(captA[23]), .A1(A[23]), .S(n20), .Z(n109) );
  CMX2X1 U949 ( .A0(captA[22]), .A1(A[22]), .S(n840), .Z(n108) );
  CMX2X1 U950 ( .A0(captA[21]), .A1(A[21]), .S(n841), .Z(n107) );
  CMX2X1 U951 ( .A0(captA[20]), .A1(A[20]), .S(n20), .Z(n106) );
  CMX2X1 U952 ( .A0(captA[19]), .A1(A[19]), .S(n840), .Z(n105) );
  CMX2X1 U953 ( .A0(captA[18]), .A1(A[18]), .S(n841), .Z(n104) );
  CMX2X1 U954 ( .A0(captA[17]), .A1(A[17]), .S(n20), .Z(n103) );
  CMX2X1 U955 ( .A0(captA[16]), .A1(A[16]), .S(n840), .Z(n102) );
  CMX2X1 U956 ( .A0(captA[15]), .A1(A[15]), .S(n841), .Z(n101) );
  CMX2X1 U957 ( .A0(captA[14]), .A1(A[14]), .S(n20), .Z(n100) );
  CMX2X1 U958 ( .A0(captA[13]), .A1(A[13]), .S(n840), .Z(n99) );
  CMX2X1 U959 ( .A0(captA[12]), .A1(A[12]), .S(n841), .Z(n98) );
  CMX2X1 U960 ( .A0(captA[11]), .A1(A[11]), .S(n20), .Z(n97) );
  CMX2X1 U961 ( .A0(captA[10]), .A1(A[10]), .S(n840), .Z(n96) );
  CMX2X1 U962 ( .A0(captA[9]), .A1(A[9]), .S(n841), .Z(n95) );
  CMX2X1 U963 ( .A0(captA[8]), .A1(A[8]), .S(n20), .Z(n94) );
  CMX2X1 U964 ( .A0(captA[7]), .A1(A[7]), .S(n840), .Z(n93) );
  CMX2X1 U965 ( .A0(captA[6]), .A1(A[6]), .S(n841), .Z(n92) );
  CMX2X1 U966 ( .A0(captA[5]), .A1(A[5]), .S(n20), .Z(n91) );
  CMX2X1 U967 ( .A0(captA[4]), .A1(A[4]), .S(n840), .Z(n90) );
  CMX2X1 U968 ( .A0(captA[3]), .A1(A[3]), .S(n841), .Z(n89) );
  CMX2X1 U969 ( .A0(captA[2]), .A1(A[2]), .S(n20), .Z(n88) );
  CMX2X1 U970 ( .A0(captA[1]), .A1(A[1]), .S(n840), .Z(n87) );
  CMX2X1 U971 ( .A0(captA[0]), .A1(A[0]), .S(n841), .Z(n86) );
  CMX2X1 U972 ( .A0(n560), .A1(B[31]), .S(n842), .Z(n85) );
  CMX2X1 U973 ( .A0(n559), .A1(B[30]), .S(n843), .Z(n84) );
  CMX2X1 U974 ( .A0(captB[29]), .A1(B[29]), .S(n18), .Z(n83) );
  CMX2X1 U975 ( .A0(n558), .A1(B[28]), .S(n842), .Z(n82) );
  CMX2X1 U976 ( .A0(captB[27]), .A1(B[27]), .S(n843), .Z(n81) );
  CMX2X1 U977 ( .A0(captB[26]), .A1(B[26]), .S(n18), .Z(n80) );
  CMX2X1 U978 ( .A0(captB[25]), .A1(B[25]), .S(n842), .Z(n79) );
  CMX2X1 U979 ( .A0(captB[24]), .A1(B[24]), .S(n843), .Z(n78) );
  CMX2X1 U980 ( .A0(captB[23]), .A1(B[23]), .S(n18), .Z(n77) );
  CMX2X1 U981 ( .A0(captB[22]), .A1(B[22]), .S(n842), .Z(n76) );
  CMX2X1 U982 ( .A0(captB[21]), .A1(B[21]), .S(n843), .Z(n75) );
  CMX2X1 U983 ( .A0(captB[20]), .A1(B[20]), .S(n18), .Z(n74) );
  CMX2X1 U984 ( .A0(captB[19]), .A1(B[19]), .S(n842), .Z(n73) );
  CMX2X1 U985 ( .A0(captB[18]), .A1(B[18]), .S(n843), .Z(n72) );
  CMX2X1 U986 ( .A0(captB[17]), .A1(B[17]), .S(n18), .Z(n71) );
  CMX2X1 U987 ( .A0(captB[16]), .A1(B[16]), .S(n842), .Z(n70) );
  CMX2X1 U988 ( .A0(captB[15]), .A1(B[15]), .S(n843), .Z(n69) );
  CMX2X1 U989 ( .A0(captB[14]), .A1(B[14]), .S(n18), .Z(n68) );
  CMX2X1 U990 ( .A0(captB[13]), .A1(B[13]), .S(n842), .Z(n67) );
  CMX2X1 U991 ( .A0(captB[12]), .A1(B[12]), .S(n843), .Z(n66) );
  CMX2X1 U992 ( .A0(captB[11]), .A1(B[11]), .S(n18), .Z(n65) );
  CMX2X1 U993 ( .A0(captB[10]), .A1(B[10]), .S(n842), .Z(n64) );
  CMX2X1 U994 ( .A0(captB[9]), .A1(B[9]), .S(n843), .Z(n63) );
  CMX2X1 U995 ( .A0(captB[8]), .A1(B[8]), .S(n18), .Z(n62) );
  CMX2X1 U996 ( .A0(captB[7]), .A1(B[7]), .S(n842), .Z(n61) );
  CMX2X1 U997 ( .A0(captB[6]), .A1(B[6]), .S(n843), .Z(n60) );
  CMX2X1 U998 ( .A0(captB[5]), .A1(B[5]), .S(n18), .Z(n59) );
  CMX2X1 U999 ( .A0(captB[4]), .A1(B[4]), .S(n842), .Z(n58) );
  CMX2X1 U1000 ( .A0(captB[3]), .A1(B[3]), .S(n843), .Z(n57) );
  CMX2X1 U1001 ( .A0(captB[2]), .A1(B[2]), .S(n18), .Z(n56) );
  CMX2X1 U1002 ( .A0(captB[1]), .A1(B[1]), .S(n842), .Z(n55) );
  CMX2X1 U1003 ( .A0(captB[0]), .A1(B[0]), .S(n843), .Z(n54) );
  CMX2X1 U1004 ( .A0(n557), .A1(C[31]), .S(n844), .Z(n53) );
  CMX2X1 U1005 ( .A0(n556), .A1(C[30]), .S(n845), .Z(n52) );
  CMX2X1 U1006 ( .A0(n555), .A1(C[29]), .S(n16), .Z(n51) );
  CMX2X1 U1007 ( .A0(n554), .A1(C[28]), .S(n844), .Z(n50) );
  CMX2X1 U1008 ( .A0(n553), .A1(C[27]), .S(n845), .Z(n49) );
  CMX2X1 U1009 ( .A0(captC[26]), .A1(C[26]), .S(n16), .Z(n48) );
  CMX2X1 U1010 ( .A0(n671), .A1(C[25]), .S(n844), .Z(n47) );
  CMX2X1 U1011 ( .A0(captC[24]), .A1(C[24]), .S(n845), .Z(n46) );
  CMX2X1 U1012 ( .A0(captC[23]), .A1(C[23]), .S(n16), .Z(n45) );
  CMX2X1 U1013 ( .A0(captC[22]), .A1(C[22]), .S(n844), .Z(n44) );
  CMX2X1 U1014 ( .A0(captC[21]), .A1(C[21]), .S(n845), .Z(n43) );
  CMX2X1 U1015 ( .A0(captC[20]), .A1(C[20]), .S(n16), .Z(n42) );
  CMX2X1 U1016 ( .A0(captC[19]), .A1(C[19]), .S(n844), .Z(n41) );
  CMX2X1 U1017 ( .A0(captC[18]), .A1(C[18]), .S(n845), .Z(n40) );
  CMX2X1 U1018 ( .A0(captC[17]), .A1(C[17]), .S(n16), .Z(n39) );
  CMX2X1 U1019 ( .A0(captC[16]), .A1(C[16]), .S(n844), .Z(n38) );
  CMX2X1 U1020 ( .A0(captC[15]), .A1(C[15]), .S(n845), .Z(n37) );
  CMX2X1 U1021 ( .A0(captC[14]), .A1(C[14]), .S(n16), .Z(n36) );
  CMX2X1 U1022 ( .A0(captC[13]), .A1(C[13]), .S(n844), .Z(n35) );
  CMX2X1 U1023 ( .A0(captC[12]), .A1(C[12]), .S(n845), .Z(n34) );
  CMX2X1 U1024 ( .A0(captC[11]), .A1(C[11]), .S(n16), .Z(n33) );
  CMX2X1 U1025 ( .A0(captC[10]), .A1(C[10]), .S(n844), .Z(n32) );
  CMX2X1 U1026 ( .A0(captC[9]), .A1(C[9]), .S(n845), .Z(n31) );
  CMX2X1 U1027 ( .A0(captC[8]), .A1(C[8]), .S(n16), .Z(n30) );
  CMX2X1 U1028 ( .A0(captC[7]), .A1(C[7]), .S(n844), .Z(n29) );
  CMX2X1 U1029 ( .A0(captC[6]), .A1(C[6]), .S(n845), .Z(n28) );
  CMX2X1 U1030 ( .A0(captC[5]), .A1(C[5]), .S(n16), .Z(n27) );
  CMX2X1 U1031 ( .A0(captC[4]), .A1(C[4]), .S(n844), .Z(n26) );
  CMX2X1 U1032 ( .A0(captC[3]), .A1(C[3]), .S(n845), .Z(n25) );
  CMX2X1 U1033 ( .A0(captC[2]), .A1(C[2]), .S(n16), .Z(n24) );
  CMX2X1 U1034 ( .A0(captC[1]), .A1(C[1]), .S(n844), .Z(n23) );
  CMX2X1 U1035 ( .A0(captC[0]), .A1(C[0]), .S(n845), .Z(n22) );
endmodule

